// -------------------------------------------------------------
//
// Module: bandpass_filter
// -------------------------------------------------------------
// HDL Implementation    : Fully parallel
// Folding Factor        : 1
// -------------------------------------------------------------



`timescale 1 ns / 1 ns

module bandpass_filter
               (
                clk,
                clk_enable,
                reset,
                filter_in,
                filter_out
                );

  input   clk; 
  input   clk_enable; 
  input   reset; 
  input   signed [15:0] filter_in; //sfix16_En15
  output  signed [35:0] filter_out; //sfix36_En34

////////////////////////////////////////////////////////////////
//Module Architecture: filter1
////////////////////////////////////////////////////////////////
  // Local Functions
  // Type Definitions
  // Constants
  parameter signed [15:0] coeff1 = 16'b0000000111010110; //sfix16_En19
  parameter signed [15:0] coeff2 = 16'b1111111111011111; //sfix16_En19
  parameter signed [15:0] coeff3 = 16'b1111111111000011; //sfix16_En19
  parameter signed [15:0] coeff4 = 16'b1111111110010101; //sfix16_En19
  parameter signed [15:0] coeff5 = 16'b1111111101010111; //sfix16_En19
  parameter signed [15:0] coeff6 = 16'b1111111100001110; //sfix16_En19
  parameter signed [15:0] coeff7 = 16'b1111111010111101; //sfix16_En19
  parameter signed [15:0] coeff8 = 16'b1111111001101010; //sfix16_En19
  parameter signed [15:0] coeff9 = 16'b1111111000011001; //sfix16_En19
  parameter signed [15:0] coeff10 = 16'b1111110111010011; //sfix16_En19
  parameter signed [15:0] coeff11 = 16'b1111110110011110; //sfix16_En19
  parameter signed [15:0] coeff12 = 16'b1111110110000000; //sfix16_En19
  parameter signed [15:0] coeff13 = 16'b1111110101111110; //sfix16_En19
  parameter signed [15:0] coeff14 = 16'b1111110110011111; //sfix16_En19
  parameter signed [15:0] coeff15 = 16'b1111110111100100; //sfix16_En19
  parameter signed [15:0] coeff16 = 16'b1111111001001111; //sfix16_En19
  parameter signed [15:0] coeff17 = 16'b1111111011011111; //sfix16_En19
  parameter signed [15:0] coeff18 = 16'b1111111110010001; //sfix16_En19
  parameter signed [15:0] coeff19 = 16'b0000000001011110; //sfix16_En19
  parameter signed [15:0] coeff20 = 16'b0000000100111111; //sfix16_En19
  parameter signed [15:0] coeff21 = 16'b0000001000101001; //sfix16_En19
  parameter signed [15:0] coeff22 = 16'b0000001100010001; //sfix16_En19
  parameter signed [15:0] coeff23 = 16'b0000001111101011; //sfix16_En19
  parameter signed [15:0] coeff24 = 16'b0000010010101010; //sfix16_En19
  parameter signed [15:0] coeff25 = 16'b0000010101000010; //sfix16_En19
  parameter signed [15:0] coeff26 = 16'b0000010110101000; //sfix16_En19
  parameter signed [15:0] coeff27 = 16'b0000010111010100; //sfix16_En19
  parameter signed [15:0] coeff28 = 16'b0000010111000001; //sfix16_En19
  parameter signed [15:0] coeff29 = 16'b0000010101101101; //sfix16_En19
  parameter signed [15:0] coeff30 = 16'b0000010011011000; //sfix16_En19
  parameter signed [15:0] coeff31 = 16'b0000010000001010; //sfix16_En19
  parameter signed [15:0] coeff32 = 16'b0000001100001011; //sfix16_En19
  parameter signed [15:0] coeff33 = 16'b0000000111100111; //sfix16_En19
  parameter signed [15:0] coeff34 = 16'b0000000010101101; //sfix16_En19
  parameter signed [15:0] coeff35 = 16'b1111111101101111; //sfix16_En19
  parameter signed [15:0] coeff36 = 16'b1111111000111110; //sfix16_En19
  parameter signed [15:0] coeff37 = 16'b1111110100101010; //sfix16_En19
  parameter signed [15:0] coeff38 = 16'b1111110001000100; //sfix16_En19
  parameter signed [15:0] coeff39 = 16'b1111101110011001; //sfix16_En19
  parameter signed [15:0] coeff40 = 16'b1111101100101111; //sfix16_En19
  parameter signed [15:0] coeff41 = 16'b1111101100001110; //sfix16_En19
  parameter signed [15:0] coeff42 = 16'b1111101100110010; //sfix16_En19
  parameter signed [15:0] coeff43 = 16'b1111101110010111; //sfix16_En19
  parameter signed [15:0] coeff44 = 16'b1111110000110000; //sfix16_En19
  parameter signed [15:0] coeff45 = 16'b1111110011101110; //sfix16_En19
  parameter signed [15:0] coeff46 = 16'b1111110110111110; //sfix16_En19
  parameter signed [15:0] coeff47 = 16'b1111111010001001; //sfix16_En19
  parameter signed [15:0] coeff48 = 16'b1111111100111001; //sfix16_En19
  parameter signed [15:0] coeff49 = 16'b1111111110111001; //sfix16_En19
  parameter signed [15:0] coeff50 = 16'b1111111111110110; //sfix16_En19
  parameter signed [15:0] coeff51 = 16'b1111111111100001; //sfix16_En19
  parameter signed [15:0] coeff52 = 16'b1111111101110001; //sfix16_En19
  parameter signed [15:0] coeff53 = 16'b1111111010100110; //sfix16_En19
  parameter signed [15:0] coeff54 = 16'b1111110110000101; //sfix16_En19
  parameter signed [15:0] coeff55 = 16'b1111110000011111; //sfix16_En19
  parameter signed [15:0] coeff56 = 16'b1111101010001000; //sfix16_En19
  parameter signed [15:0] coeff57 = 16'b1111100011100000; //sfix16_En19
  parameter signed [15:0] coeff58 = 16'b1111011101001010; //sfix16_En19
  parameter signed [15:0] coeff59 = 16'b1111010111101101; //sfix16_En19
  parameter signed [15:0] coeff60 = 16'b1111010011110010; //sfix16_En19
  parameter signed [15:0] coeff61 = 16'b1111010010000000; //sfix16_En19
  parameter signed [15:0] coeff62 = 16'b1111010010111011; //sfix16_En19
  parameter signed [15:0] coeff63 = 16'b1111010110111101; //sfix16_En19
  parameter signed [15:0] coeff64 = 16'b1111011110011001; //sfix16_En19
  parameter signed [15:0] coeff65 = 16'b1111101001010110; //sfix16_En19
  parameter signed [15:0] coeff66 = 16'b1111110111101100; //sfix16_En19
  parameter signed [15:0] coeff67 = 16'b0000001001000100; //sfix16_En19
  parameter signed [15:0] coeff68 = 16'b0000011100111011; //sfix16_En19
  parameter signed [15:0] coeff69 = 16'b0000110010011110; //sfix16_En19
  parameter signed [15:0] coeff70 = 16'b0001001000101110; //sfix16_En19
  parameter signed [15:0] coeff71 = 16'b0001011110100100; //sfix16_En19
  parameter signed [15:0] coeff72 = 16'b0001110010110000; //sfix16_En19
  parameter signed [15:0] coeff73 = 16'b0010000100000100; //sfix16_En19
  parameter signed [15:0] coeff74 = 16'b0010010001001111; //sfix16_En19
  parameter signed [15:0] coeff75 = 16'b0010011001001100; //sfix16_En19
  parameter signed [15:0] coeff76 = 16'b0010011010111111; //sfix16_En19
  parameter signed [15:0] coeff77 = 16'b0010010101111010; //sfix16_En19
  parameter signed [15:0] coeff78 = 16'b0010001001100110; //sfix16_En19
  parameter signed [15:0] coeff79 = 16'b0001110110000000; //sfix16_En19
  parameter signed [15:0] coeff80 = 16'b0001011011011100; //sfix16_En19
  parameter signed [15:0] coeff81 = 16'b0000111010100111; //sfix16_En19
  parameter signed [15:0] coeff82 = 16'b0000010100100110; //sfix16_En19
  parameter signed [15:0] coeff83 = 16'b1111101010110010; //sfix16_En19
  parameter signed [15:0] coeff84 = 16'b1110111110110110; //sfix16_En19
  parameter signed [15:0] coeff85 = 16'b1110010010101100; //sfix16_En19
  parameter signed [15:0] coeff86 = 16'b1101101000010011; //sfix16_En19
  parameter signed [15:0] coeff87 = 16'b1101000001101111; //sfix16_En19
  parameter signed [15:0] coeff88 = 16'b1100100000111011; //sfix16_En19
  parameter signed [15:0] coeff89 = 16'b1100000111101011; //sfix16_En19
  parameter signed [15:0] coeff90 = 16'b1011110111011101; //sfix16_En19
  parameter signed [15:0] coeff91 = 16'b1011110001011101; //sfix16_En19
  parameter signed [15:0] coeff92 = 16'b1011110110010101; //sfix16_En19
  parameter signed [15:0] coeff93 = 16'b1100000110010110; //sfix16_En19
  parameter signed [15:0] coeff94 = 16'b1100100001001101; //sfix16_En19
  parameter signed [15:0] coeff95 = 16'b1101000110000111; //sfix16_En19
  parameter signed [15:0] coeff96 = 16'b1101110011110001; //sfix16_En19
  parameter signed [15:0] coeff97 = 16'b1110101000011100; //sfix16_En19
  parameter signed [15:0] coeff98 = 16'b1111100010000011; //sfix16_En19
  parameter signed [15:0] coeff99 = 16'b0000011110001101; //sfix16_En19
  parameter signed [15:0] coeff100 = 16'b0001011010011001; //sfix16_En19
  parameter signed [15:0] coeff101 = 16'b0010010100000000; //sfix16_En19
  parameter signed [15:0] coeff102 = 16'b0011001000100010; //sfix16_En19
  parameter signed [15:0] coeff103 = 16'b0011110101101011; //sfix16_En19
  parameter signed [15:0] coeff104 = 16'b0100011001011011; //sfix16_En19
  parameter signed [15:0] coeff105 = 16'b0100110010001100; //sfix16_En19
  parameter signed [15:0] coeff106 = 16'b0100111110110111; //sfix16_En19
  parameter signed [15:0] coeff107 = 16'b0100111110110111; //sfix16_En19
  parameter signed [15:0] coeff108 = 16'b0100110010001100; //sfix16_En19
  parameter signed [15:0] coeff109 = 16'b0100011001011011; //sfix16_En19
  parameter signed [15:0] coeff110 = 16'b0011110101101011; //sfix16_En19
  parameter signed [15:0] coeff111 = 16'b0011001000100010; //sfix16_En19
  parameter signed [15:0] coeff112 = 16'b0010010100000000; //sfix16_En19
  parameter signed [15:0] coeff113 = 16'b0001011010011001; //sfix16_En19
  parameter signed [15:0] coeff114 = 16'b0000011110001101; //sfix16_En19
  parameter signed [15:0] coeff115 = 16'b1111100010000011; //sfix16_En19
  parameter signed [15:0] coeff116 = 16'b1110101000011100; //sfix16_En19
  parameter signed [15:0] coeff117 = 16'b1101110011110001; //sfix16_En19
  parameter signed [15:0] coeff118 = 16'b1101000110000111; //sfix16_En19
  parameter signed [15:0] coeff119 = 16'b1100100001001101; //sfix16_En19
  parameter signed [15:0] coeff120 = 16'b1100000110010110; //sfix16_En19
  parameter signed [15:0] coeff121 = 16'b1011110110010101; //sfix16_En19
  parameter signed [15:0] coeff122 = 16'b1011110001011101; //sfix16_En19
  parameter signed [15:0] coeff123 = 16'b1011110111011101; //sfix16_En19
  parameter signed [15:0] coeff124 = 16'b1100000111101011; //sfix16_En19
  parameter signed [15:0] coeff125 = 16'b1100100000111011; //sfix16_En19
  parameter signed [15:0] coeff126 = 16'b1101000001101111; //sfix16_En19
  parameter signed [15:0] coeff127 = 16'b1101101000010011; //sfix16_En19
  parameter signed [15:0] coeff128 = 16'b1110010010101100; //sfix16_En19
  parameter signed [15:0] coeff129 = 16'b1110111110110110; //sfix16_En19
  parameter signed [15:0] coeff130 = 16'b1111101010110010; //sfix16_En19
  parameter signed [15:0] coeff131 = 16'b0000010100100110; //sfix16_En19
  parameter signed [15:0] coeff132 = 16'b0000111010100111; //sfix16_En19
  parameter signed [15:0] coeff133 = 16'b0001011011011100; //sfix16_En19
  parameter signed [15:0] coeff134 = 16'b0001110110000000; //sfix16_En19
  parameter signed [15:0] coeff135 = 16'b0010001001100110; //sfix16_En19
  parameter signed [15:0] coeff136 = 16'b0010010101111010; //sfix16_En19
  parameter signed [15:0] coeff137 = 16'b0010011010111111; //sfix16_En19
  parameter signed [15:0] coeff138 = 16'b0010011001001100; //sfix16_En19
  parameter signed [15:0] coeff139 = 16'b0010010001001111; //sfix16_En19
  parameter signed [15:0] coeff140 = 16'b0010000100000100; //sfix16_En19
  parameter signed [15:0] coeff141 = 16'b0001110010110000; //sfix16_En19
  parameter signed [15:0] coeff142 = 16'b0001011110100100; //sfix16_En19
  parameter signed [15:0] coeff143 = 16'b0001001000101110; //sfix16_En19
  parameter signed [15:0] coeff144 = 16'b0000110010011110; //sfix16_En19
  parameter signed [15:0] coeff145 = 16'b0000011100111011; //sfix16_En19
  parameter signed [15:0] coeff146 = 16'b0000001001000100; //sfix16_En19
  parameter signed [15:0] coeff147 = 16'b1111110111101100; //sfix16_En19
  parameter signed [15:0] coeff148 = 16'b1111101001010110; //sfix16_En19
  parameter signed [15:0] coeff149 = 16'b1111011110011001; //sfix16_En19
  parameter signed [15:0] coeff150 = 16'b1111010110111101; //sfix16_En19
  parameter signed [15:0] coeff151 = 16'b1111010010111011; //sfix16_En19
  parameter signed [15:0] coeff152 = 16'b1111010010000000; //sfix16_En19
  parameter signed [15:0] coeff153 = 16'b1111010011110010; //sfix16_En19
  parameter signed [15:0] coeff154 = 16'b1111010111101101; //sfix16_En19
  parameter signed [15:0] coeff155 = 16'b1111011101001010; //sfix16_En19
  parameter signed [15:0] coeff156 = 16'b1111100011100000; //sfix16_En19
  parameter signed [15:0] coeff157 = 16'b1111101010001000; //sfix16_En19
  parameter signed [15:0] coeff158 = 16'b1111110000011111; //sfix16_En19
  parameter signed [15:0] coeff159 = 16'b1111110110000101; //sfix16_En19
  parameter signed [15:0] coeff160 = 16'b1111111010100110; //sfix16_En19
  parameter signed [15:0] coeff161 = 16'b1111111101110001; //sfix16_En19
  parameter signed [15:0] coeff162 = 16'b1111111111100001; //sfix16_En19
  parameter signed [15:0] coeff163 = 16'b1111111111110110; //sfix16_En19
  parameter signed [15:0] coeff164 = 16'b1111111110111001; //sfix16_En19
  parameter signed [15:0] coeff165 = 16'b1111111100111001; //sfix16_En19
  parameter signed [15:0] coeff166 = 16'b1111111010001001; //sfix16_En19
  parameter signed [15:0] coeff167 = 16'b1111110110111110; //sfix16_En19
  parameter signed [15:0] coeff168 = 16'b1111110011101110; //sfix16_En19
  parameter signed [15:0] coeff169 = 16'b1111110000110000; //sfix16_En19
  parameter signed [15:0] coeff170 = 16'b1111101110010111; //sfix16_En19
  parameter signed [15:0] coeff171 = 16'b1111101100110010; //sfix16_En19
  parameter signed [15:0] coeff172 = 16'b1111101100001110; //sfix16_En19
  parameter signed [15:0] coeff173 = 16'b1111101100101111; //sfix16_En19
  parameter signed [15:0] coeff174 = 16'b1111101110011001; //sfix16_En19
  parameter signed [15:0] coeff175 = 16'b1111110001000100; //sfix16_En19
  parameter signed [15:0] coeff176 = 16'b1111110100101010; //sfix16_En19
  parameter signed [15:0] coeff177 = 16'b1111111000111110; //sfix16_En19
  parameter signed [15:0] coeff178 = 16'b1111111101101111; //sfix16_En19
  parameter signed [15:0] coeff179 = 16'b0000000010101101; //sfix16_En19
  parameter signed [15:0] coeff180 = 16'b0000000111100111; //sfix16_En19
  parameter signed [15:0] coeff181 = 16'b0000001100001011; //sfix16_En19
  parameter signed [15:0] coeff182 = 16'b0000010000001010; //sfix16_En19
  parameter signed [15:0] coeff183 = 16'b0000010011011000; //sfix16_En19
  parameter signed [15:0] coeff184 = 16'b0000010101101101; //sfix16_En19
  parameter signed [15:0] coeff185 = 16'b0000010111000001; //sfix16_En19
  parameter signed [15:0] coeff186 = 16'b0000010111010100; //sfix16_En19
  parameter signed [15:0] coeff187 = 16'b0000010110101000; //sfix16_En19
  parameter signed [15:0] coeff188 = 16'b0000010101000010; //sfix16_En19
  parameter signed [15:0] coeff189 = 16'b0000010010101010; //sfix16_En19
  parameter signed [15:0] coeff190 = 16'b0000001111101011; //sfix16_En19
  parameter signed [15:0] coeff191 = 16'b0000001100010001; //sfix16_En19
  parameter signed [15:0] coeff192 = 16'b0000001000101001; //sfix16_En19
  parameter signed [15:0] coeff193 = 16'b0000000100111111; //sfix16_En19
  parameter signed [15:0] coeff194 = 16'b0000000001011110; //sfix16_En19
  parameter signed [15:0] coeff195 = 16'b1111111110010001; //sfix16_En19
  parameter signed [15:0] coeff196 = 16'b1111111011011111; //sfix16_En19
  parameter signed [15:0] coeff197 = 16'b1111111001001111; //sfix16_En19
  parameter signed [15:0] coeff198 = 16'b1111110111100100; //sfix16_En19
  parameter signed [15:0] coeff199 = 16'b1111110110011111; //sfix16_En19
  parameter signed [15:0] coeff200 = 16'b1111110101111110; //sfix16_En19
  parameter signed [15:0] coeff201 = 16'b1111110110000000; //sfix16_En19
  parameter signed [15:0] coeff202 = 16'b1111110110011110; //sfix16_En19
  parameter signed [15:0] coeff203 = 16'b1111110111010011; //sfix16_En19
  parameter signed [15:0] coeff204 = 16'b1111111000011001; //sfix16_En19
  parameter signed [15:0] coeff205 = 16'b1111111001101010; //sfix16_En19
  parameter signed [15:0] coeff206 = 16'b1111111010111101; //sfix16_En19
  parameter signed [15:0] coeff207 = 16'b1111111100001110; //sfix16_En19
  parameter signed [15:0] coeff208 = 16'b1111111101010111; //sfix16_En19
  parameter signed [15:0] coeff209 = 16'b1111111110010101; //sfix16_En19
  parameter signed [15:0] coeff210 = 16'b1111111111000011; //sfix16_En19
  parameter signed [15:0] coeff211 = 16'b1111111111011111; //sfix16_En19
  parameter signed [15:0] coeff212 = 16'b0000000111010110; //sfix16_En19

  // Signals
  reg  signed [15:0] delay_pipeline [0:211] ; // sfix16_En15
  wire signed [30:0] product212; // sfix31_En34
  wire signed [31:0] mul_temp; // sfix32_En34
  wire signed [30:0] product211; // sfix31_En34
  wire signed [31:0] mul_temp_1; // sfix32_En34
  wire signed [30:0] product210; // sfix31_En34
  wire signed [31:0] mul_temp_2; // sfix32_En34
  wire signed [30:0] product209; // sfix31_En34
  wire signed [31:0] mul_temp_3; // sfix32_En34
  wire signed [30:0] product208; // sfix31_En34
  wire signed [31:0] mul_temp_4; // sfix32_En34
  wire signed [30:0] product207; // sfix31_En34
  wire signed [31:0] mul_temp_5; // sfix32_En34
  wire signed [30:0] product206; // sfix31_En34
  wire signed [31:0] mul_temp_6; // sfix32_En34
  wire signed [30:0] product205; // sfix31_En34
  wire signed [31:0] mul_temp_7; // sfix32_En34
  wire signed [30:0] product204; // sfix31_En34
  wire signed [31:0] mul_temp_8; // sfix32_En34
  wire signed [30:0] product203; // sfix31_En34
  wire signed [31:0] mul_temp_9; // sfix32_En34
  wire signed [30:0] product202; // sfix31_En34
  wire signed [31:0] mul_temp_10; // sfix32_En34
  wire signed [30:0] product201; // sfix31_En34
  wire signed [31:0] mul_temp_11; // sfix32_En34
  wire signed [30:0] product200; // sfix31_En34
  wire signed [31:0] mul_temp_12; // sfix32_En34
  wire signed [30:0] product199; // sfix31_En34
  wire signed [31:0] mul_temp_13; // sfix32_En34
  wire signed [30:0] product198; // sfix31_En34
  wire signed [31:0] mul_temp_14; // sfix32_En34
  wire signed [30:0] product197; // sfix31_En34
  wire signed [31:0] mul_temp_15; // sfix32_En34
  wire signed [30:0] product196; // sfix31_En34
  wire signed [31:0] mul_temp_16; // sfix32_En34
  wire signed [30:0] product195; // sfix31_En34
  wire signed [31:0] mul_temp_17; // sfix32_En34
  wire signed [30:0] product194; // sfix31_En34
  wire signed [31:0] mul_temp_18; // sfix32_En34
  wire signed [30:0] product193; // sfix31_En34
  wire signed [31:0] mul_temp_19; // sfix32_En34
  wire signed [30:0] product192; // sfix31_En34
  wire signed [31:0] mul_temp_20; // sfix32_En34
  wire signed [30:0] product191; // sfix31_En34
  wire signed [31:0] mul_temp_21; // sfix32_En34
  wire signed [30:0] product190; // sfix31_En34
  wire signed [31:0] mul_temp_22; // sfix32_En34
  wire signed [30:0] product189; // sfix31_En34
  wire signed [31:0] mul_temp_23; // sfix32_En34
  wire signed [30:0] product188; // sfix31_En34
  wire signed [31:0] mul_temp_24; // sfix32_En34
  wire signed [30:0] product187; // sfix31_En34
  wire signed [31:0] mul_temp_25; // sfix32_En34
  wire signed [30:0] product186; // sfix31_En34
  wire signed [31:0] mul_temp_26; // sfix32_En34
  wire signed [30:0] product185; // sfix31_En34
  wire signed [31:0] mul_temp_27; // sfix32_En34
  wire signed [30:0] product184; // sfix31_En34
  wire signed [31:0] mul_temp_28; // sfix32_En34
  wire signed [30:0] product183; // sfix31_En34
  wire signed [31:0] mul_temp_29; // sfix32_En34
  wire signed [30:0] product182; // sfix31_En34
  wire signed [31:0] mul_temp_30; // sfix32_En34
  wire signed [30:0] product181; // sfix31_En34
  wire signed [31:0] mul_temp_31; // sfix32_En34
  wire signed [30:0] product180; // sfix31_En34
  wire signed [31:0] mul_temp_32; // sfix32_En34
  wire signed [30:0] product179; // sfix31_En34
  wire signed [31:0] mul_temp_33; // sfix32_En34
  wire signed [30:0] product178; // sfix31_En34
  wire signed [31:0] mul_temp_34; // sfix32_En34
  wire signed [30:0] product177; // sfix31_En34
  wire signed [31:0] mul_temp_35; // sfix32_En34
  wire signed [30:0] product176; // sfix31_En34
  wire signed [31:0] mul_temp_36; // sfix32_En34
  wire signed [30:0] product175; // sfix31_En34
  wire signed [31:0] mul_temp_37; // sfix32_En34
  wire signed [30:0] product174; // sfix31_En34
  wire signed [31:0] mul_temp_38; // sfix32_En34
  wire signed [30:0] product173; // sfix31_En34
  wire signed [31:0] mul_temp_39; // sfix32_En34
  wire signed [30:0] product172; // sfix31_En34
  wire signed [31:0] mul_temp_40; // sfix32_En34
  wire signed [30:0] product171; // sfix31_En34
  wire signed [31:0] mul_temp_41; // sfix32_En34
  wire signed [30:0] product170; // sfix31_En34
  wire signed [31:0] mul_temp_42; // sfix32_En34
  wire signed [30:0] product169; // sfix31_En34
  wire signed [31:0] mul_temp_43; // sfix32_En34
  wire signed [30:0] product168; // sfix31_En34
  wire signed [31:0] mul_temp_44; // sfix32_En34
  wire signed [30:0] product167; // sfix31_En34
  wire signed [31:0] mul_temp_45; // sfix32_En34
  wire signed [30:0] product166; // sfix31_En34
  wire signed [31:0] mul_temp_46; // sfix32_En34
  wire signed [30:0] product165; // sfix31_En34
  wire signed [31:0] mul_temp_47; // sfix32_En34
  wire signed [30:0] product164; // sfix31_En34
  wire signed [31:0] mul_temp_48; // sfix32_En34
  wire signed [30:0] product163; // sfix31_En34
  wire signed [31:0] mul_temp_49; // sfix32_En34
  wire signed [30:0] product162; // sfix31_En34
  wire signed [31:0] mul_temp_50; // sfix32_En34
  wire signed [30:0] product161; // sfix31_En34
  wire signed [31:0] mul_temp_51; // sfix32_En34
  wire signed [30:0] product160; // sfix31_En34
  wire signed [31:0] mul_temp_52; // sfix32_En34
  wire signed [30:0] product159; // sfix31_En34
  wire signed [31:0] mul_temp_53; // sfix32_En34
  wire signed [30:0] product158; // sfix31_En34
  wire signed [31:0] mul_temp_54; // sfix32_En34
  wire signed [30:0] product157; // sfix31_En34
  wire signed [31:0] mul_temp_55; // sfix32_En34
  wire signed [30:0] product156; // sfix31_En34
  wire signed [31:0] mul_temp_56; // sfix32_En34
  wire signed [30:0] product155; // sfix31_En34
  wire signed [31:0] mul_temp_57; // sfix32_En34
  wire signed [30:0] product154; // sfix31_En34
  wire signed [31:0] mul_temp_58; // sfix32_En34
  wire signed [30:0] product153; // sfix31_En34
  wire signed [31:0] mul_temp_59; // sfix32_En34
  wire signed [30:0] product152; // sfix31_En34
  wire signed [31:0] mul_temp_60; // sfix32_En34
  wire signed [30:0] product151; // sfix31_En34
  wire signed [31:0] mul_temp_61; // sfix32_En34
  wire signed [30:0] product150; // sfix31_En34
  wire signed [31:0] mul_temp_62; // sfix32_En34
  wire signed [30:0] product149; // sfix31_En34
  wire signed [31:0] mul_temp_63; // sfix32_En34
  wire signed [30:0] product148; // sfix31_En34
  wire signed [31:0] mul_temp_64; // sfix32_En34
  wire signed [30:0] product147; // sfix31_En34
  wire signed [31:0] mul_temp_65; // sfix32_En34
  wire signed [30:0] product146; // sfix31_En34
  wire signed [31:0] mul_temp_66; // sfix32_En34
  wire signed [30:0] product145; // sfix31_En34
  wire signed [31:0] mul_temp_67; // sfix32_En34
  wire signed [30:0] product144; // sfix31_En34
  wire signed [31:0] mul_temp_68; // sfix32_En34
  wire signed [30:0] product143; // sfix31_En34
  wire signed [31:0] mul_temp_69; // sfix32_En34
  wire signed [30:0] product142; // sfix31_En34
  wire signed [31:0] mul_temp_70; // sfix32_En34
  wire signed [30:0] product141; // sfix31_En34
  wire signed [31:0] mul_temp_71; // sfix32_En34
  wire signed [30:0] product140; // sfix31_En34
  wire signed [31:0] mul_temp_72; // sfix32_En34
  wire signed [30:0] product139; // sfix31_En34
  wire signed [31:0] mul_temp_73; // sfix32_En34
  wire signed [30:0] product138; // sfix31_En34
  wire signed [31:0] mul_temp_74; // sfix32_En34
  wire signed [30:0] product137; // sfix31_En34
  wire signed [31:0] mul_temp_75; // sfix32_En34
  wire signed [30:0] product136; // sfix31_En34
  wire signed [31:0] mul_temp_76; // sfix32_En34
  wire signed [30:0] product135; // sfix31_En34
  wire signed [31:0] mul_temp_77; // sfix32_En34
  wire signed [30:0] product134; // sfix31_En34
  wire signed [31:0] mul_temp_78; // sfix32_En34
  wire signed [30:0] product133; // sfix31_En34
  wire signed [31:0] mul_temp_79; // sfix32_En34
  wire signed [30:0] product132; // sfix31_En34
  wire signed [31:0] mul_temp_80; // sfix32_En34
  wire signed [30:0] product131; // sfix31_En34
  wire signed [31:0] mul_temp_81; // sfix32_En34
  wire signed [30:0] product130; // sfix31_En34
  wire signed [31:0] mul_temp_82; // sfix32_En34
  wire signed [30:0] product129; // sfix31_En34
  wire signed [31:0] mul_temp_83; // sfix32_En34
  wire signed [30:0] product128; // sfix31_En34
  wire signed [31:0] mul_temp_84; // sfix32_En34
  wire signed [30:0] product127; // sfix31_En34
  wire signed [31:0] mul_temp_85; // sfix32_En34
  wire signed [30:0] product126; // sfix31_En34
  wire signed [31:0] mul_temp_86; // sfix32_En34
  wire signed [30:0] product125; // sfix31_En34
  wire signed [31:0] mul_temp_87; // sfix32_En34
  wire signed [30:0] product124; // sfix31_En34
  wire signed [31:0] mul_temp_88; // sfix32_En34
  wire signed [30:0] product123; // sfix31_En34
  wire signed [31:0] mul_temp_89; // sfix32_En34
  wire signed [30:0] product122; // sfix31_En34
  wire signed [31:0] mul_temp_90; // sfix32_En34
  wire signed [30:0] product121; // sfix31_En34
  wire signed [31:0] mul_temp_91; // sfix32_En34
  wire signed [30:0] product120; // sfix31_En34
  wire signed [31:0] mul_temp_92; // sfix32_En34
  wire signed [30:0] product119; // sfix31_En34
  wire signed [31:0] mul_temp_93; // sfix32_En34
  wire signed [30:0] product118; // sfix31_En34
  wire signed [31:0] mul_temp_94; // sfix32_En34
  wire signed [30:0] product117; // sfix31_En34
  wire signed [31:0] mul_temp_95; // sfix32_En34
  wire signed [30:0] product116; // sfix31_En34
  wire signed [31:0] mul_temp_96; // sfix32_En34
  wire signed [30:0] product115; // sfix31_En34
  wire signed [31:0] mul_temp_97; // sfix32_En34
  wire signed [30:0] product114; // sfix31_En34
  wire signed [31:0] mul_temp_98; // sfix32_En34
  wire signed [30:0] product113; // sfix31_En34
  wire signed [31:0] mul_temp_99; // sfix32_En34
  wire signed [30:0] product112; // sfix31_En34
  wire signed [31:0] mul_temp_100; // sfix32_En34
  wire signed [30:0] product111; // sfix31_En34
  wire signed [31:0] mul_temp_101; // sfix32_En34
  wire signed [30:0] product110; // sfix31_En34
  wire signed [31:0] mul_temp_102; // sfix32_En34
  wire signed [30:0] product109; // sfix31_En34
  wire signed [31:0] mul_temp_103; // sfix32_En34
  wire signed [30:0] product108; // sfix31_En34
  wire signed [31:0] mul_temp_104; // sfix32_En34
  wire signed [30:0] product107; // sfix31_En34
  wire signed [31:0] mul_temp_105; // sfix32_En34
  wire signed [30:0] product106; // sfix31_En34
  wire signed [31:0] mul_temp_106; // sfix32_En34
  wire signed [30:0] product105; // sfix31_En34
  wire signed [31:0] mul_temp_107; // sfix32_En34
  wire signed [30:0] product104; // sfix31_En34
  wire signed [31:0] mul_temp_108; // sfix32_En34
  wire signed [30:0] product103; // sfix31_En34
  wire signed [31:0] mul_temp_109; // sfix32_En34
  wire signed [30:0] product102; // sfix31_En34
  wire signed [31:0] mul_temp_110; // sfix32_En34
  wire signed [30:0] product101; // sfix31_En34
  wire signed [31:0] mul_temp_111; // sfix32_En34
  wire signed [30:0] product100; // sfix31_En34
  wire signed [31:0] mul_temp_112; // sfix32_En34
  wire signed [30:0] product99; // sfix31_En34
  wire signed [31:0] mul_temp_113; // sfix32_En34
  wire signed [30:0] product98; // sfix31_En34
  wire signed [31:0] mul_temp_114; // sfix32_En34
  wire signed [30:0] product97; // sfix31_En34
  wire signed [31:0] mul_temp_115; // sfix32_En34
  wire signed [30:0] product96; // sfix31_En34
  wire signed [31:0] mul_temp_116; // sfix32_En34
  wire signed [30:0] product95; // sfix31_En34
  wire signed [31:0] mul_temp_117; // sfix32_En34
  wire signed [30:0] product94; // sfix31_En34
  wire signed [31:0] mul_temp_118; // sfix32_En34
  wire signed [30:0] product93; // sfix31_En34
  wire signed [31:0] mul_temp_119; // sfix32_En34
  wire signed [30:0] product92; // sfix31_En34
  wire signed [31:0] mul_temp_120; // sfix32_En34
  wire signed [30:0] product91; // sfix31_En34
  wire signed [31:0] mul_temp_121; // sfix32_En34
  wire signed [30:0] product90; // sfix31_En34
  wire signed [31:0] mul_temp_122; // sfix32_En34
  wire signed [30:0] product89; // sfix31_En34
  wire signed [31:0] mul_temp_123; // sfix32_En34
  wire signed [30:0] product88; // sfix31_En34
  wire signed [31:0] mul_temp_124; // sfix32_En34
  wire signed [30:0] product87; // sfix31_En34
  wire signed [31:0] mul_temp_125; // sfix32_En34
  wire signed [30:0] product86; // sfix31_En34
  wire signed [31:0] mul_temp_126; // sfix32_En34
  wire signed [30:0] product85; // sfix31_En34
  wire signed [31:0] mul_temp_127; // sfix32_En34
  wire signed [30:0] product84; // sfix31_En34
  wire signed [31:0] mul_temp_128; // sfix32_En34
  wire signed [30:0] product83; // sfix31_En34
  wire signed [31:0] mul_temp_129; // sfix32_En34
  wire signed [30:0] product82; // sfix31_En34
  wire signed [31:0] mul_temp_130; // sfix32_En34
  wire signed [30:0] product81; // sfix31_En34
  wire signed [31:0] mul_temp_131; // sfix32_En34
  wire signed [30:0] product80; // sfix31_En34
  wire signed [31:0] mul_temp_132; // sfix32_En34
  wire signed [30:0] product79; // sfix31_En34
  wire signed [31:0] mul_temp_133; // sfix32_En34
  wire signed [30:0] product78; // sfix31_En34
  wire signed [31:0] mul_temp_134; // sfix32_En34
  wire signed [30:0] product77; // sfix31_En34
  wire signed [31:0] mul_temp_135; // sfix32_En34
  wire signed [30:0] product76; // sfix31_En34
  wire signed [31:0] mul_temp_136; // sfix32_En34
  wire signed [30:0] product75; // sfix31_En34
  wire signed [31:0] mul_temp_137; // sfix32_En34
  wire signed [30:0] product74; // sfix31_En34
  wire signed [31:0] mul_temp_138; // sfix32_En34
  wire signed [30:0] product73; // sfix31_En34
  wire signed [31:0] mul_temp_139; // sfix32_En34
  wire signed [30:0] product72; // sfix31_En34
  wire signed [31:0] mul_temp_140; // sfix32_En34
  wire signed [30:0] product71; // sfix31_En34
  wire signed [31:0] mul_temp_141; // sfix32_En34
  wire signed [30:0] product70; // sfix31_En34
  wire signed [31:0] mul_temp_142; // sfix32_En34
  wire signed [30:0] product69; // sfix31_En34
  wire signed [31:0] mul_temp_143; // sfix32_En34
  wire signed [30:0] product68; // sfix31_En34
  wire signed [31:0] mul_temp_144; // sfix32_En34
  wire signed [30:0] product67; // sfix31_En34
  wire signed [31:0] mul_temp_145; // sfix32_En34
  wire signed [30:0] product66; // sfix31_En34
  wire signed [31:0] mul_temp_146; // sfix32_En34
  wire signed [30:0] product65; // sfix31_En34
  wire signed [31:0] mul_temp_147; // sfix32_En34
  wire signed [30:0] product64; // sfix31_En34
  wire signed [31:0] mul_temp_148; // sfix32_En34
  wire signed [30:0] product63; // sfix31_En34
  wire signed [31:0] mul_temp_149; // sfix32_En34
  wire signed [30:0] product62; // sfix31_En34
  wire signed [31:0] mul_temp_150; // sfix32_En34
  wire signed [30:0] product61; // sfix31_En34
  wire signed [31:0] mul_temp_151; // sfix32_En34
  wire signed [30:0] product60; // sfix31_En34
  wire signed [31:0] mul_temp_152; // sfix32_En34
  wire signed [30:0] product59; // sfix31_En34
  wire signed [31:0] mul_temp_153; // sfix32_En34
  wire signed [30:0] product58; // sfix31_En34
  wire signed [31:0] mul_temp_154; // sfix32_En34
  wire signed [30:0] product57; // sfix31_En34
  wire signed [31:0] mul_temp_155; // sfix32_En34
  wire signed [30:0] product56; // sfix31_En34
  wire signed [31:0] mul_temp_156; // sfix32_En34
  wire signed [30:0] product55; // sfix31_En34
  wire signed [31:0] mul_temp_157; // sfix32_En34
  wire signed [30:0] product54; // sfix31_En34
  wire signed [31:0] mul_temp_158; // sfix32_En34
  wire signed [30:0] product53; // sfix31_En34
  wire signed [31:0] mul_temp_159; // sfix32_En34
  wire signed [30:0] product52; // sfix31_En34
  wire signed [31:0] mul_temp_160; // sfix32_En34
  wire signed [30:0] product51; // sfix31_En34
  wire signed [31:0] mul_temp_161; // sfix32_En34
  wire signed [30:0] product50; // sfix31_En34
  wire signed [31:0] mul_temp_162; // sfix32_En34
  wire signed [30:0] product49; // sfix31_En34
  wire signed [31:0] mul_temp_163; // sfix32_En34
  wire signed [30:0] product48; // sfix31_En34
  wire signed [31:0] mul_temp_164; // sfix32_En34
  wire signed [30:0] product47; // sfix31_En34
  wire signed [31:0] mul_temp_165; // sfix32_En34
  wire signed [30:0] product46; // sfix31_En34
  wire signed [31:0] mul_temp_166; // sfix32_En34
  wire signed [30:0] product45; // sfix31_En34
  wire signed [31:0] mul_temp_167; // sfix32_En34
  wire signed [30:0] product44; // sfix31_En34
  wire signed [31:0] mul_temp_168; // sfix32_En34
  wire signed [30:0] product43; // sfix31_En34
  wire signed [31:0] mul_temp_169; // sfix32_En34
  wire signed [30:0] product42; // sfix31_En34
  wire signed [31:0] mul_temp_170; // sfix32_En34
  wire signed [30:0] product41; // sfix31_En34
  wire signed [31:0] mul_temp_171; // sfix32_En34
  wire signed [30:0] product40; // sfix31_En34
  wire signed [31:0] mul_temp_172; // sfix32_En34
  wire signed [30:0] product39; // sfix31_En34
  wire signed [31:0] mul_temp_173; // sfix32_En34
  wire signed [30:0] product38; // sfix31_En34
  wire signed [31:0] mul_temp_174; // sfix32_En34
  wire signed [30:0] product37; // sfix31_En34
  wire signed [31:0] mul_temp_175; // sfix32_En34
  wire signed [30:0] product36; // sfix31_En34
  wire signed [31:0] mul_temp_176; // sfix32_En34
  wire signed [30:0] product35; // sfix31_En34
  wire signed [31:0] mul_temp_177; // sfix32_En34
  wire signed [30:0] product34; // sfix31_En34
  wire signed [31:0] mul_temp_178; // sfix32_En34
  wire signed [30:0] product33; // sfix31_En34
  wire signed [31:0] mul_temp_179; // sfix32_En34
  wire signed [30:0] product32; // sfix31_En34
  wire signed [31:0] mul_temp_180; // sfix32_En34
  wire signed [30:0] product31; // sfix31_En34
  wire signed [31:0] mul_temp_181; // sfix32_En34
  wire signed [30:0] product30; // sfix31_En34
  wire signed [31:0] mul_temp_182; // sfix32_En34
  wire signed [30:0] product29; // sfix31_En34
  wire signed [31:0] mul_temp_183; // sfix32_En34
  wire signed [30:0] product28; // sfix31_En34
  wire signed [31:0] mul_temp_184; // sfix32_En34
  wire signed [30:0] product27; // sfix31_En34
  wire signed [31:0] mul_temp_185; // sfix32_En34
  wire signed [30:0] product26; // sfix31_En34
  wire signed [31:0] mul_temp_186; // sfix32_En34
  wire signed [30:0] product25; // sfix31_En34
  wire signed [31:0] mul_temp_187; // sfix32_En34
  wire signed [30:0] product24; // sfix31_En34
  wire signed [31:0] mul_temp_188; // sfix32_En34
  wire signed [30:0] product23; // sfix31_En34
  wire signed [31:0] mul_temp_189; // sfix32_En34
  wire signed [30:0] product22; // sfix31_En34
  wire signed [31:0] mul_temp_190; // sfix32_En34
  wire signed [30:0] product21; // sfix31_En34
  wire signed [31:0] mul_temp_191; // sfix32_En34
  wire signed [30:0] product20; // sfix31_En34
  wire signed [31:0] mul_temp_192; // sfix32_En34
  wire signed [30:0] product19; // sfix31_En34
  wire signed [31:0] mul_temp_193; // sfix32_En34
  wire signed [30:0] product18; // sfix31_En34
  wire signed [31:0] mul_temp_194; // sfix32_En34
  wire signed [30:0] product17; // sfix31_En34
  wire signed [31:0] mul_temp_195; // sfix32_En34
  wire signed [30:0] product16; // sfix31_En34
  wire signed [31:0] mul_temp_196; // sfix32_En34
  wire signed [30:0] product15; // sfix31_En34
  wire signed [31:0] mul_temp_197; // sfix32_En34
  wire signed [30:0] product14; // sfix31_En34
  wire signed [31:0] mul_temp_198; // sfix32_En34
  wire signed [30:0] product13; // sfix31_En34
  wire signed [31:0] mul_temp_199; // sfix32_En34
  wire signed [30:0] product12; // sfix31_En34
  wire signed [31:0] mul_temp_200; // sfix32_En34
  wire signed [30:0] product11; // sfix31_En34
  wire signed [31:0] mul_temp_201; // sfix32_En34
  wire signed [30:0] product10; // sfix31_En34
  wire signed [31:0] mul_temp_202; // sfix32_En34
  wire signed [30:0] product9; // sfix31_En34
  wire signed [31:0] mul_temp_203; // sfix32_En34
  wire signed [30:0] product8; // sfix31_En34
  wire signed [31:0] mul_temp_204; // sfix32_En34
  wire signed [30:0] product7; // sfix31_En34
  wire signed [31:0] mul_temp_205; // sfix32_En34
  wire signed [30:0] product6; // sfix31_En34
  wire signed [31:0] mul_temp_206; // sfix32_En34
  wire signed [30:0] product5; // sfix31_En34
  wire signed [31:0] mul_temp_207; // sfix32_En34
  wire signed [30:0] product4; // sfix31_En34
  wire signed [31:0] mul_temp_208; // sfix32_En34
  wire signed [30:0] product3; // sfix31_En34
  wire signed [31:0] mul_temp_209; // sfix32_En34
  wire signed [30:0] product2; // sfix31_En34
  wire signed [31:0] mul_temp_210; // sfix32_En34
  wire signed [35:0] product1_cast; // sfix36_En34
  wire signed [30:0] product1; // sfix31_En34
  wire signed [31:0] mul_temp_211; // sfix32_En34
  wire signed [35:0] sum1; // sfix36_En34
  wire signed [35:0] add_signext; // sfix36_En34
  wire signed [35:0] add_signext_1; // sfix36_En34
  wire signed [36:0] add_temp; // sfix37_En34
  wire signed [35:0] sum2; // sfix36_En34
  wire signed [35:0] add_signext_2; // sfix36_En34
  wire signed [35:0] add_signext_3; // sfix36_En34
  wire signed [36:0] add_temp_1; // sfix37_En34
  wire signed [35:0] sum3; // sfix36_En34
  wire signed [35:0] add_signext_4; // sfix36_En34
  wire signed [35:0] add_signext_5; // sfix36_En34
  wire signed [36:0] add_temp_2; // sfix37_En34
  wire signed [35:0] sum4; // sfix36_En34
  wire signed [35:0] add_signext_6; // sfix36_En34
  wire signed [35:0] add_signext_7; // sfix36_En34
  wire signed [36:0] add_temp_3; // sfix37_En34
  wire signed [35:0] sum5; // sfix36_En34
  wire signed [35:0] add_signext_8; // sfix36_En34
  wire signed [35:0] add_signext_9; // sfix36_En34
  wire signed [36:0] add_temp_4; // sfix37_En34
  wire signed [35:0] sum6; // sfix36_En34
  wire signed [35:0] add_signext_10; // sfix36_En34
  wire signed [35:0] add_signext_11; // sfix36_En34
  wire signed [36:0] add_temp_5; // sfix37_En34
  wire signed [35:0] sum7; // sfix36_En34
  wire signed [35:0] add_signext_12; // sfix36_En34
  wire signed [35:0] add_signext_13; // sfix36_En34
  wire signed [36:0] add_temp_6; // sfix37_En34
  wire signed [35:0] sum8; // sfix36_En34
  wire signed [35:0] add_signext_14; // sfix36_En34
  wire signed [35:0] add_signext_15; // sfix36_En34
  wire signed [36:0] add_temp_7; // sfix37_En34
  wire signed [35:0] sum9; // sfix36_En34
  wire signed [35:0] add_signext_16; // sfix36_En34
  wire signed [35:0] add_signext_17; // sfix36_En34
  wire signed [36:0] add_temp_8; // sfix37_En34
  wire signed [35:0] sum10; // sfix36_En34
  wire signed [35:0] add_signext_18; // sfix36_En34
  wire signed [35:0] add_signext_19; // sfix36_En34
  wire signed [36:0] add_temp_9; // sfix37_En34
  wire signed [35:0] sum11; // sfix36_En34
  wire signed [35:0] add_signext_20; // sfix36_En34
  wire signed [35:0] add_signext_21; // sfix36_En34
  wire signed [36:0] add_temp_10; // sfix37_En34
  wire signed [35:0] sum12; // sfix36_En34
  wire signed [35:0] add_signext_22; // sfix36_En34
  wire signed [35:0] add_signext_23; // sfix36_En34
  wire signed [36:0] add_temp_11; // sfix37_En34
  wire signed [35:0] sum13; // sfix36_En34
  wire signed [35:0] add_signext_24; // sfix36_En34
  wire signed [35:0] add_signext_25; // sfix36_En34
  wire signed [36:0] add_temp_12; // sfix37_En34
  wire signed [35:0] sum14; // sfix36_En34
  wire signed [35:0] add_signext_26; // sfix36_En34
  wire signed [35:0] add_signext_27; // sfix36_En34
  wire signed [36:0] add_temp_13; // sfix37_En34
  wire signed [35:0] sum15; // sfix36_En34
  wire signed [35:0] add_signext_28; // sfix36_En34
  wire signed [35:0] add_signext_29; // sfix36_En34
  wire signed [36:0] add_temp_14; // sfix37_En34
  wire signed [35:0] sum16; // sfix36_En34
  wire signed [35:0] add_signext_30; // sfix36_En34
  wire signed [35:0] add_signext_31; // sfix36_En34
  wire signed [36:0] add_temp_15; // sfix37_En34
  wire signed [35:0] sum17; // sfix36_En34
  wire signed [35:0] add_signext_32; // sfix36_En34
  wire signed [35:0] add_signext_33; // sfix36_En34
  wire signed [36:0] add_temp_16; // sfix37_En34
  wire signed [35:0] sum18; // sfix36_En34
  wire signed [35:0] add_signext_34; // sfix36_En34
  wire signed [35:0] add_signext_35; // sfix36_En34
  wire signed [36:0] add_temp_17; // sfix37_En34
  wire signed [35:0] sum19; // sfix36_En34
  wire signed [35:0] add_signext_36; // sfix36_En34
  wire signed [35:0] add_signext_37; // sfix36_En34
  wire signed [36:0] add_temp_18; // sfix37_En34
  wire signed [35:0] sum20; // sfix36_En34
  wire signed [35:0] add_signext_38; // sfix36_En34
  wire signed [35:0] add_signext_39; // sfix36_En34
  wire signed [36:0] add_temp_19; // sfix37_En34
  wire signed [35:0] sum21; // sfix36_En34
  wire signed [35:0] add_signext_40; // sfix36_En34
  wire signed [35:0] add_signext_41; // sfix36_En34
  wire signed [36:0] add_temp_20; // sfix37_En34
  wire signed [35:0] sum22; // sfix36_En34
  wire signed [35:0] add_signext_42; // sfix36_En34
  wire signed [35:0] add_signext_43; // sfix36_En34
  wire signed [36:0] add_temp_21; // sfix37_En34
  wire signed [35:0] sum23; // sfix36_En34
  wire signed [35:0] add_signext_44; // sfix36_En34
  wire signed [35:0] add_signext_45; // sfix36_En34
  wire signed [36:0] add_temp_22; // sfix37_En34
  wire signed [35:0] sum24; // sfix36_En34
  wire signed [35:0] add_signext_46; // sfix36_En34
  wire signed [35:0] add_signext_47; // sfix36_En34
  wire signed [36:0] add_temp_23; // sfix37_En34
  wire signed [35:0] sum25; // sfix36_En34
  wire signed [35:0] add_signext_48; // sfix36_En34
  wire signed [35:0] add_signext_49; // sfix36_En34
  wire signed [36:0] add_temp_24; // sfix37_En34
  wire signed [35:0] sum26; // sfix36_En34
  wire signed [35:0] add_signext_50; // sfix36_En34
  wire signed [35:0] add_signext_51; // sfix36_En34
  wire signed [36:0] add_temp_25; // sfix37_En34
  wire signed [35:0] sum27; // sfix36_En34
  wire signed [35:0] add_signext_52; // sfix36_En34
  wire signed [35:0] add_signext_53; // sfix36_En34
  wire signed [36:0] add_temp_26; // sfix37_En34
  wire signed [35:0] sum28; // sfix36_En34
  wire signed [35:0] add_signext_54; // sfix36_En34
  wire signed [35:0] add_signext_55; // sfix36_En34
  wire signed [36:0] add_temp_27; // sfix37_En34
  wire signed [35:0] sum29; // sfix36_En34
  wire signed [35:0] add_signext_56; // sfix36_En34
  wire signed [35:0] add_signext_57; // sfix36_En34
  wire signed [36:0] add_temp_28; // sfix37_En34
  wire signed [35:0] sum30; // sfix36_En34
  wire signed [35:0] add_signext_58; // sfix36_En34
  wire signed [35:0] add_signext_59; // sfix36_En34
  wire signed [36:0] add_temp_29; // sfix37_En34
  wire signed [35:0] sum31; // sfix36_En34
  wire signed [35:0] add_signext_60; // sfix36_En34
  wire signed [35:0] add_signext_61; // sfix36_En34
  wire signed [36:0] add_temp_30; // sfix37_En34
  wire signed [35:0] sum32; // sfix36_En34
  wire signed [35:0] add_signext_62; // sfix36_En34
  wire signed [35:0] add_signext_63; // sfix36_En34
  wire signed [36:0] add_temp_31; // sfix37_En34
  wire signed [35:0] sum33; // sfix36_En34
  wire signed [35:0] add_signext_64; // sfix36_En34
  wire signed [35:0] add_signext_65; // sfix36_En34
  wire signed [36:0] add_temp_32; // sfix37_En34
  wire signed [35:0] sum34; // sfix36_En34
  wire signed [35:0] add_signext_66; // sfix36_En34
  wire signed [35:0] add_signext_67; // sfix36_En34
  wire signed [36:0] add_temp_33; // sfix37_En34
  wire signed [35:0] sum35; // sfix36_En34
  wire signed [35:0] add_signext_68; // sfix36_En34
  wire signed [35:0] add_signext_69; // sfix36_En34
  wire signed [36:0] add_temp_34; // sfix37_En34
  wire signed [35:0] sum36; // sfix36_En34
  wire signed [35:0] add_signext_70; // sfix36_En34
  wire signed [35:0] add_signext_71; // sfix36_En34
  wire signed [36:0] add_temp_35; // sfix37_En34
  wire signed [35:0] sum37; // sfix36_En34
  wire signed [35:0] add_signext_72; // sfix36_En34
  wire signed [35:0] add_signext_73; // sfix36_En34
  wire signed [36:0] add_temp_36; // sfix37_En34
  wire signed [35:0] sum38; // sfix36_En34
  wire signed [35:0] add_signext_74; // sfix36_En34
  wire signed [35:0] add_signext_75; // sfix36_En34
  wire signed [36:0] add_temp_37; // sfix37_En34
  wire signed [35:0] sum39; // sfix36_En34
  wire signed [35:0] add_signext_76; // sfix36_En34
  wire signed [35:0] add_signext_77; // sfix36_En34
  wire signed [36:0] add_temp_38; // sfix37_En34
  wire signed [35:0] sum40; // sfix36_En34
  wire signed [35:0] add_signext_78; // sfix36_En34
  wire signed [35:0] add_signext_79; // sfix36_En34
  wire signed [36:0] add_temp_39; // sfix37_En34
  wire signed [35:0] sum41; // sfix36_En34
  wire signed [35:0] add_signext_80; // sfix36_En34
  wire signed [35:0] add_signext_81; // sfix36_En34
  wire signed [36:0] add_temp_40; // sfix37_En34
  wire signed [35:0] sum42; // sfix36_En34
  wire signed [35:0] add_signext_82; // sfix36_En34
  wire signed [35:0] add_signext_83; // sfix36_En34
  wire signed [36:0] add_temp_41; // sfix37_En34
  wire signed [35:0] sum43; // sfix36_En34
  wire signed [35:0] add_signext_84; // sfix36_En34
  wire signed [35:0] add_signext_85; // sfix36_En34
  wire signed [36:0] add_temp_42; // sfix37_En34
  wire signed [35:0] sum44; // sfix36_En34
  wire signed [35:0] add_signext_86; // sfix36_En34
  wire signed [35:0] add_signext_87; // sfix36_En34
  wire signed [36:0] add_temp_43; // sfix37_En34
  wire signed [35:0] sum45; // sfix36_En34
  wire signed [35:0] add_signext_88; // sfix36_En34
  wire signed [35:0] add_signext_89; // sfix36_En34
  wire signed [36:0] add_temp_44; // sfix37_En34
  wire signed [35:0] sum46; // sfix36_En34
  wire signed [35:0] add_signext_90; // sfix36_En34
  wire signed [35:0] add_signext_91; // sfix36_En34
  wire signed [36:0] add_temp_45; // sfix37_En34
  wire signed [35:0] sum47; // sfix36_En34
  wire signed [35:0] add_signext_92; // sfix36_En34
  wire signed [35:0] add_signext_93; // sfix36_En34
  wire signed [36:0] add_temp_46; // sfix37_En34
  wire signed [35:0] sum48; // sfix36_En34
  wire signed [35:0] add_signext_94; // sfix36_En34
  wire signed [35:0] add_signext_95; // sfix36_En34
  wire signed [36:0] add_temp_47; // sfix37_En34
  wire signed [35:0] sum49; // sfix36_En34
  wire signed [35:0] add_signext_96; // sfix36_En34
  wire signed [35:0] add_signext_97; // sfix36_En34
  wire signed [36:0] add_temp_48; // sfix37_En34
  wire signed [35:0] sum50; // sfix36_En34
  wire signed [35:0] add_signext_98; // sfix36_En34
  wire signed [35:0] add_signext_99; // sfix36_En34
  wire signed [36:0] add_temp_49; // sfix37_En34
  wire signed [35:0] sum51; // sfix36_En34
  wire signed [35:0] add_signext_100; // sfix36_En34
  wire signed [35:0] add_signext_101; // sfix36_En34
  wire signed [36:0] add_temp_50; // sfix37_En34
  wire signed [35:0] sum52; // sfix36_En34
  wire signed [35:0] add_signext_102; // sfix36_En34
  wire signed [35:0] add_signext_103; // sfix36_En34
  wire signed [36:0] add_temp_51; // sfix37_En34
  wire signed [35:0] sum53; // sfix36_En34
  wire signed [35:0] add_signext_104; // sfix36_En34
  wire signed [35:0] add_signext_105; // sfix36_En34
  wire signed [36:0] add_temp_52; // sfix37_En34
  wire signed [35:0] sum54; // sfix36_En34
  wire signed [35:0] add_signext_106; // sfix36_En34
  wire signed [35:0] add_signext_107; // sfix36_En34
  wire signed [36:0] add_temp_53; // sfix37_En34
  wire signed [35:0] sum55; // sfix36_En34
  wire signed [35:0] add_signext_108; // sfix36_En34
  wire signed [35:0] add_signext_109; // sfix36_En34
  wire signed [36:0] add_temp_54; // sfix37_En34
  wire signed [35:0] sum56; // sfix36_En34
  wire signed [35:0] add_signext_110; // sfix36_En34
  wire signed [35:0] add_signext_111; // sfix36_En34
  wire signed [36:0] add_temp_55; // sfix37_En34
  wire signed [35:0] sum57; // sfix36_En34
  wire signed [35:0] add_signext_112; // sfix36_En34
  wire signed [35:0] add_signext_113; // sfix36_En34
  wire signed [36:0] add_temp_56; // sfix37_En34
  wire signed [35:0] sum58; // sfix36_En34
  wire signed [35:0] add_signext_114; // sfix36_En34
  wire signed [35:0] add_signext_115; // sfix36_En34
  wire signed [36:0] add_temp_57; // sfix37_En34
  wire signed [35:0] sum59; // sfix36_En34
  wire signed [35:0] add_signext_116; // sfix36_En34
  wire signed [35:0] add_signext_117; // sfix36_En34
  wire signed [36:0] add_temp_58; // sfix37_En34
  wire signed [35:0] sum60; // sfix36_En34
  wire signed [35:0] add_signext_118; // sfix36_En34
  wire signed [35:0] add_signext_119; // sfix36_En34
  wire signed [36:0] add_temp_59; // sfix37_En34
  wire signed [35:0] sum61; // sfix36_En34
  wire signed [35:0] add_signext_120; // sfix36_En34
  wire signed [35:0] add_signext_121; // sfix36_En34
  wire signed [36:0] add_temp_60; // sfix37_En34
  wire signed [35:0] sum62; // sfix36_En34
  wire signed [35:0] add_signext_122; // sfix36_En34
  wire signed [35:0] add_signext_123; // sfix36_En34
  wire signed [36:0] add_temp_61; // sfix37_En34
  wire signed [35:0] sum63; // sfix36_En34
  wire signed [35:0] add_signext_124; // sfix36_En34
  wire signed [35:0] add_signext_125; // sfix36_En34
  wire signed [36:0] add_temp_62; // sfix37_En34
  wire signed [35:0] sum64; // sfix36_En34
  wire signed [35:0] add_signext_126; // sfix36_En34
  wire signed [35:0] add_signext_127; // sfix36_En34
  wire signed [36:0] add_temp_63; // sfix37_En34
  wire signed [35:0] sum65; // sfix36_En34
  wire signed [35:0] add_signext_128; // sfix36_En34
  wire signed [35:0] add_signext_129; // sfix36_En34
  wire signed [36:0] add_temp_64; // sfix37_En34
  wire signed [35:0] sum66; // sfix36_En34
  wire signed [35:0] add_signext_130; // sfix36_En34
  wire signed [35:0] add_signext_131; // sfix36_En34
  wire signed [36:0] add_temp_65; // sfix37_En34
  wire signed [35:0] sum67; // sfix36_En34
  wire signed [35:0] add_signext_132; // sfix36_En34
  wire signed [35:0] add_signext_133; // sfix36_En34
  wire signed [36:0] add_temp_66; // sfix37_En34
  wire signed [35:0] sum68; // sfix36_En34
  wire signed [35:0] add_signext_134; // sfix36_En34
  wire signed [35:0] add_signext_135; // sfix36_En34
  wire signed [36:0] add_temp_67; // sfix37_En34
  wire signed [35:0] sum69; // sfix36_En34
  wire signed [35:0] add_signext_136; // sfix36_En34
  wire signed [35:0] add_signext_137; // sfix36_En34
  wire signed [36:0] add_temp_68; // sfix37_En34
  wire signed [35:0] sum70; // sfix36_En34
  wire signed [35:0] add_signext_138; // sfix36_En34
  wire signed [35:0] add_signext_139; // sfix36_En34
  wire signed [36:0] add_temp_69; // sfix37_En34
  wire signed [35:0] sum71; // sfix36_En34
  wire signed [35:0] add_signext_140; // sfix36_En34
  wire signed [35:0] add_signext_141; // sfix36_En34
  wire signed [36:0] add_temp_70; // sfix37_En34
  wire signed [35:0] sum72; // sfix36_En34
  wire signed [35:0] add_signext_142; // sfix36_En34
  wire signed [35:0] add_signext_143; // sfix36_En34
  wire signed [36:0] add_temp_71; // sfix37_En34
  wire signed [35:0] sum73; // sfix36_En34
  wire signed [35:0] add_signext_144; // sfix36_En34
  wire signed [35:0] add_signext_145; // sfix36_En34
  wire signed [36:0] add_temp_72; // sfix37_En34
  wire signed [35:0] sum74; // sfix36_En34
  wire signed [35:0] add_signext_146; // sfix36_En34
  wire signed [35:0] add_signext_147; // sfix36_En34
  wire signed [36:0] add_temp_73; // sfix37_En34
  wire signed [35:0] sum75; // sfix36_En34
  wire signed [35:0] add_signext_148; // sfix36_En34
  wire signed [35:0] add_signext_149; // sfix36_En34
  wire signed [36:0] add_temp_74; // sfix37_En34
  wire signed [35:0] sum76; // sfix36_En34
  wire signed [35:0] add_signext_150; // sfix36_En34
  wire signed [35:0] add_signext_151; // sfix36_En34
  wire signed [36:0] add_temp_75; // sfix37_En34
  wire signed [35:0] sum77; // sfix36_En34
  wire signed [35:0] add_signext_152; // sfix36_En34
  wire signed [35:0] add_signext_153; // sfix36_En34
  wire signed [36:0] add_temp_76; // sfix37_En34
  wire signed [35:0] sum78; // sfix36_En34
  wire signed [35:0] add_signext_154; // sfix36_En34
  wire signed [35:0] add_signext_155; // sfix36_En34
  wire signed [36:0] add_temp_77; // sfix37_En34
  wire signed [35:0] sum79; // sfix36_En34
  wire signed [35:0] add_signext_156; // sfix36_En34
  wire signed [35:0] add_signext_157; // sfix36_En34
  wire signed [36:0] add_temp_78; // sfix37_En34
  wire signed [35:0] sum80; // sfix36_En34
  wire signed [35:0] add_signext_158; // sfix36_En34
  wire signed [35:0] add_signext_159; // sfix36_En34
  wire signed [36:0] add_temp_79; // sfix37_En34
  wire signed [35:0] sum81; // sfix36_En34
  wire signed [35:0] add_signext_160; // sfix36_En34
  wire signed [35:0] add_signext_161; // sfix36_En34
  wire signed [36:0] add_temp_80; // sfix37_En34
  wire signed [35:0] sum82; // sfix36_En34
  wire signed [35:0] add_signext_162; // sfix36_En34
  wire signed [35:0] add_signext_163; // sfix36_En34
  wire signed [36:0] add_temp_81; // sfix37_En34
  wire signed [35:0] sum83; // sfix36_En34
  wire signed [35:0] add_signext_164; // sfix36_En34
  wire signed [35:0] add_signext_165; // sfix36_En34
  wire signed [36:0] add_temp_82; // sfix37_En34
  wire signed [35:0] sum84; // sfix36_En34
  wire signed [35:0] add_signext_166; // sfix36_En34
  wire signed [35:0] add_signext_167; // sfix36_En34
  wire signed [36:0] add_temp_83; // sfix37_En34
  wire signed [35:0] sum85; // sfix36_En34
  wire signed [35:0] add_signext_168; // sfix36_En34
  wire signed [35:0] add_signext_169; // sfix36_En34
  wire signed [36:0] add_temp_84; // sfix37_En34
  wire signed [35:0] sum86; // sfix36_En34
  wire signed [35:0] add_signext_170; // sfix36_En34
  wire signed [35:0] add_signext_171; // sfix36_En34
  wire signed [36:0] add_temp_85; // sfix37_En34
  wire signed [35:0] sum87; // sfix36_En34
  wire signed [35:0] add_signext_172; // sfix36_En34
  wire signed [35:0] add_signext_173; // sfix36_En34
  wire signed [36:0] add_temp_86; // sfix37_En34
  wire signed [35:0] sum88; // sfix36_En34
  wire signed [35:0] add_signext_174; // sfix36_En34
  wire signed [35:0] add_signext_175; // sfix36_En34
  wire signed [36:0] add_temp_87; // sfix37_En34
  wire signed [35:0] sum89; // sfix36_En34
  wire signed [35:0] add_signext_176; // sfix36_En34
  wire signed [35:0] add_signext_177; // sfix36_En34
  wire signed [36:0] add_temp_88; // sfix37_En34
  wire signed [35:0] sum90; // sfix36_En34
  wire signed [35:0] add_signext_178; // sfix36_En34
  wire signed [35:0] add_signext_179; // sfix36_En34
  wire signed [36:0] add_temp_89; // sfix37_En34
  wire signed [35:0] sum91; // sfix36_En34
  wire signed [35:0] add_signext_180; // sfix36_En34
  wire signed [35:0] add_signext_181; // sfix36_En34
  wire signed [36:0] add_temp_90; // sfix37_En34
  wire signed [35:0] sum92; // sfix36_En34
  wire signed [35:0] add_signext_182; // sfix36_En34
  wire signed [35:0] add_signext_183; // sfix36_En34
  wire signed [36:0] add_temp_91; // sfix37_En34
  wire signed [35:0] sum93; // sfix36_En34
  wire signed [35:0] add_signext_184; // sfix36_En34
  wire signed [35:0] add_signext_185; // sfix36_En34
  wire signed [36:0] add_temp_92; // sfix37_En34
  wire signed [35:0] sum94; // sfix36_En34
  wire signed [35:0] add_signext_186; // sfix36_En34
  wire signed [35:0] add_signext_187; // sfix36_En34
  wire signed [36:0] add_temp_93; // sfix37_En34
  wire signed [35:0] sum95; // sfix36_En34
  wire signed [35:0] add_signext_188; // sfix36_En34
  wire signed [35:0] add_signext_189; // sfix36_En34
  wire signed [36:0] add_temp_94; // sfix37_En34
  wire signed [35:0] sum96; // sfix36_En34
  wire signed [35:0] add_signext_190; // sfix36_En34
  wire signed [35:0] add_signext_191; // sfix36_En34
  wire signed [36:0] add_temp_95; // sfix37_En34
  wire signed [35:0] sum97; // sfix36_En34
  wire signed [35:0] add_signext_192; // sfix36_En34
  wire signed [35:0] add_signext_193; // sfix36_En34
  wire signed [36:0] add_temp_96; // sfix37_En34
  wire signed [35:0] sum98; // sfix36_En34
  wire signed [35:0] add_signext_194; // sfix36_En34
  wire signed [35:0] add_signext_195; // sfix36_En34
  wire signed [36:0] add_temp_97; // sfix37_En34
  wire signed [35:0] sum99; // sfix36_En34
  wire signed [35:0] add_signext_196; // sfix36_En34
  wire signed [35:0] add_signext_197; // sfix36_En34
  wire signed [36:0] add_temp_98; // sfix37_En34
  wire signed [35:0] sum100; // sfix36_En34
  wire signed [35:0] add_signext_198; // sfix36_En34
  wire signed [35:0] add_signext_199; // sfix36_En34
  wire signed [36:0] add_temp_99; // sfix37_En34
  wire signed [35:0] sum101; // sfix36_En34
  wire signed [35:0] add_signext_200; // sfix36_En34
  wire signed [35:0] add_signext_201; // sfix36_En34
  wire signed [36:0] add_temp_100; // sfix37_En34
  wire signed [35:0] sum102; // sfix36_En34
  wire signed [35:0] add_signext_202; // sfix36_En34
  wire signed [35:0] add_signext_203; // sfix36_En34
  wire signed [36:0] add_temp_101; // sfix37_En34
  wire signed [35:0] sum103; // sfix36_En34
  wire signed [35:0] add_signext_204; // sfix36_En34
  wire signed [35:0] add_signext_205; // sfix36_En34
  wire signed [36:0] add_temp_102; // sfix37_En34
  wire signed [35:0] sum104; // sfix36_En34
  wire signed [35:0] add_signext_206; // sfix36_En34
  wire signed [35:0] add_signext_207; // sfix36_En34
  wire signed [36:0] add_temp_103; // sfix37_En34
  wire signed [35:0] sum105; // sfix36_En34
  wire signed [35:0] add_signext_208; // sfix36_En34
  wire signed [35:0] add_signext_209; // sfix36_En34
  wire signed [36:0] add_temp_104; // sfix37_En34
  wire signed [35:0] sum106; // sfix36_En34
  wire signed [35:0] add_signext_210; // sfix36_En34
  wire signed [35:0] add_signext_211; // sfix36_En34
  wire signed [36:0] add_temp_105; // sfix37_En34
  wire signed [35:0] sum107; // sfix36_En34
  wire signed [35:0] add_signext_212; // sfix36_En34
  wire signed [35:0] add_signext_213; // sfix36_En34
  wire signed [36:0] add_temp_106; // sfix37_En34
  wire signed [35:0] sum108; // sfix36_En34
  wire signed [35:0] add_signext_214; // sfix36_En34
  wire signed [35:0] add_signext_215; // sfix36_En34
  wire signed [36:0] add_temp_107; // sfix37_En34
  wire signed [35:0] sum109; // sfix36_En34
  wire signed [35:0] add_signext_216; // sfix36_En34
  wire signed [35:0] add_signext_217; // sfix36_En34
  wire signed [36:0] add_temp_108; // sfix37_En34
  wire signed [35:0] sum110; // sfix36_En34
  wire signed [35:0] add_signext_218; // sfix36_En34
  wire signed [35:0] add_signext_219; // sfix36_En34
  wire signed [36:0] add_temp_109; // sfix37_En34
  wire signed [35:0] sum111; // sfix36_En34
  wire signed [35:0] add_signext_220; // sfix36_En34
  wire signed [35:0] add_signext_221; // sfix36_En34
  wire signed [36:0] add_temp_110; // sfix37_En34
  wire signed [35:0] sum112; // sfix36_En34
  wire signed [35:0] add_signext_222; // sfix36_En34
  wire signed [35:0] add_signext_223; // sfix36_En34
  wire signed [36:0] add_temp_111; // sfix37_En34
  wire signed [35:0] sum113; // sfix36_En34
  wire signed [35:0] add_signext_224; // sfix36_En34
  wire signed [35:0] add_signext_225; // sfix36_En34
  wire signed [36:0] add_temp_112; // sfix37_En34
  wire signed [35:0] sum114; // sfix36_En34
  wire signed [35:0] add_signext_226; // sfix36_En34
  wire signed [35:0] add_signext_227; // sfix36_En34
  wire signed [36:0] add_temp_113; // sfix37_En34
  wire signed [35:0] sum115; // sfix36_En34
  wire signed [35:0] add_signext_228; // sfix36_En34
  wire signed [35:0] add_signext_229; // sfix36_En34
  wire signed [36:0] add_temp_114; // sfix37_En34
  wire signed [35:0] sum116; // sfix36_En34
  wire signed [35:0] add_signext_230; // sfix36_En34
  wire signed [35:0] add_signext_231; // sfix36_En34
  wire signed [36:0] add_temp_115; // sfix37_En34
  wire signed [35:0] sum117; // sfix36_En34
  wire signed [35:0] add_signext_232; // sfix36_En34
  wire signed [35:0] add_signext_233; // sfix36_En34
  wire signed [36:0] add_temp_116; // sfix37_En34
  wire signed [35:0] sum118; // sfix36_En34
  wire signed [35:0] add_signext_234; // sfix36_En34
  wire signed [35:0] add_signext_235; // sfix36_En34
  wire signed [36:0] add_temp_117; // sfix37_En34
  wire signed [35:0] sum119; // sfix36_En34
  wire signed [35:0] add_signext_236; // sfix36_En34
  wire signed [35:0] add_signext_237; // sfix36_En34
  wire signed [36:0] add_temp_118; // sfix37_En34
  wire signed [35:0] sum120; // sfix36_En34
  wire signed [35:0] add_signext_238; // sfix36_En34
  wire signed [35:0] add_signext_239; // sfix36_En34
  wire signed [36:0] add_temp_119; // sfix37_En34
  wire signed [35:0] sum121; // sfix36_En34
  wire signed [35:0] add_signext_240; // sfix36_En34
  wire signed [35:0] add_signext_241; // sfix36_En34
  wire signed [36:0] add_temp_120; // sfix37_En34
  wire signed [35:0] sum122; // sfix36_En34
  wire signed [35:0] add_signext_242; // sfix36_En34
  wire signed [35:0] add_signext_243; // sfix36_En34
  wire signed [36:0] add_temp_121; // sfix37_En34
  wire signed [35:0] sum123; // sfix36_En34
  wire signed [35:0] add_signext_244; // sfix36_En34
  wire signed [35:0] add_signext_245; // sfix36_En34
  wire signed [36:0] add_temp_122; // sfix37_En34
  wire signed [35:0] sum124; // sfix36_En34
  wire signed [35:0] add_signext_246; // sfix36_En34
  wire signed [35:0] add_signext_247; // sfix36_En34
  wire signed [36:0] add_temp_123; // sfix37_En34
  wire signed [35:0] sum125; // sfix36_En34
  wire signed [35:0] add_signext_248; // sfix36_En34
  wire signed [35:0] add_signext_249; // sfix36_En34
  wire signed [36:0] add_temp_124; // sfix37_En34
  wire signed [35:0] sum126; // sfix36_En34
  wire signed [35:0] add_signext_250; // sfix36_En34
  wire signed [35:0] add_signext_251; // sfix36_En34
  wire signed [36:0] add_temp_125; // sfix37_En34
  wire signed [35:0] sum127; // sfix36_En34
  wire signed [35:0] add_signext_252; // sfix36_En34
  wire signed [35:0] add_signext_253; // sfix36_En34
  wire signed [36:0] add_temp_126; // sfix37_En34
  wire signed [35:0] sum128; // sfix36_En34
  wire signed [35:0] add_signext_254; // sfix36_En34
  wire signed [35:0] add_signext_255; // sfix36_En34
  wire signed [36:0] add_temp_127; // sfix37_En34
  wire signed [35:0] sum129; // sfix36_En34
  wire signed [35:0] add_signext_256; // sfix36_En34
  wire signed [35:0] add_signext_257; // sfix36_En34
  wire signed [36:0] add_temp_128; // sfix37_En34
  wire signed [35:0] sum130; // sfix36_En34
  wire signed [35:0] add_signext_258; // sfix36_En34
  wire signed [35:0] add_signext_259; // sfix36_En34
  wire signed [36:0] add_temp_129; // sfix37_En34
  wire signed [35:0] sum131; // sfix36_En34
  wire signed [35:0] add_signext_260; // sfix36_En34
  wire signed [35:0] add_signext_261; // sfix36_En34
  wire signed [36:0] add_temp_130; // sfix37_En34
  wire signed [35:0] sum132; // sfix36_En34
  wire signed [35:0] add_signext_262; // sfix36_En34
  wire signed [35:0] add_signext_263; // sfix36_En34
  wire signed [36:0] add_temp_131; // sfix37_En34
  wire signed [35:0] sum133; // sfix36_En34
  wire signed [35:0] add_signext_264; // sfix36_En34
  wire signed [35:0] add_signext_265; // sfix36_En34
  wire signed [36:0] add_temp_132; // sfix37_En34
  wire signed [35:0] sum134; // sfix36_En34
  wire signed [35:0] add_signext_266; // sfix36_En34
  wire signed [35:0] add_signext_267; // sfix36_En34
  wire signed [36:0] add_temp_133; // sfix37_En34
  wire signed [35:0] sum135; // sfix36_En34
  wire signed [35:0] add_signext_268; // sfix36_En34
  wire signed [35:0] add_signext_269; // sfix36_En34
  wire signed [36:0] add_temp_134; // sfix37_En34
  wire signed [35:0] sum136; // sfix36_En34
  wire signed [35:0] add_signext_270; // sfix36_En34
  wire signed [35:0] add_signext_271; // sfix36_En34
  wire signed [36:0] add_temp_135; // sfix37_En34
  wire signed [35:0] sum137; // sfix36_En34
  wire signed [35:0] add_signext_272; // sfix36_En34
  wire signed [35:0] add_signext_273; // sfix36_En34
  wire signed [36:0] add_temp_136; // sfix37_En34
  wire signed [35:0] sum138; // sfix36_En34
  wire signed [35:0] add_signext_274; // sfix36_En34
  wire signed [35:0] add_signext_275; // sfix36_En34
  wire signed [36:0] add_temp_137; // sfix37_En34
  wire signed [35:0] sum139; // sfix36_En34
  wire signed [35:0] add_signext_276; // sfix36_En34
  wire signed [35:0] add_signext_277; // sfix36_En34
  wire signed [36:0] add_temp_138; // sfix37_En34
  wire signed [35:0] sum140; // sfix36_En34
  wire signed [35:0] add_signext_278; // sfix36_En34
  wire signed [35:0] add_signext_279; // sfix36_En34
  wire signed [36:0] add_temp_139; // sfix37_En34
  wire signed [35:0] sum141; // sfix36_En34
  wire signed [35:0] add_signext_280; // sfix36_En34
  wire signed [35:0] add_signext_281; // sfix36_En34
  wire signed [36:0] add_temp_140; // sfix37_En34
  wire signed [35:0] sum142; // sfix36_En34
  wire signed [35:0] add_signext_282; // sfix36_En34
  wire signed [35:0] add_signext_283; // sfix36_En34
  wire signed [36:0] add_temp_141; // sfix37_En34
  wire signed [35:0] sum143; // sfix36_En34
  wire signed [35:0] add_signext_284; // sfix36_En34
  wire signed [35:0] add_signext_285; // sfix36_En34
  wire signed [36:0] add_temp_142; // sfix37_En34
  wire signed [35:0] sum144; // sfix36_En34
  wire signed [35:0] add_signext_286; // sfix36_En34
  wire signed [35:0] add_signext_287; // sfix36_En34
  wire signed [36:0] add_temp_143; // sfix37_En34
  wire signed [35:0] sum145; // sfix36_En34
  wire signed [35:0] add_signext_288; // sfix36_En34
  wire signed [35:0] add_signext_289; // sfix36_En34
  wire signed [36:0] add_temp_144; // sfix37_En34
  wire signed [35:0] sum146; // sfix36_En34
  wire signed [35:0] add_signext_290; // sfix36_En34
  wire signed [35:0] add_signext_291; // sfix36_En34
  wire signed [36:0] add_temp_145; // sfix37_En34
  wire signed [35:0] sum147; // sfix36_En34
  wire signed [35:0] add_signext_292; // sfix36_En34
  wire signed [35:0] add_signext_293; // sfix36_En34
  wire signed [36:0] add_temp_146; // sfix37_En34
  wire signed [35:0] sum148; // sfix36_En34
  wire signed [35:0] add_signext_294; // sfix36_En34
  wire signed [35:0] add_signext_295; // sfix36_En34
  wire signed [36:0] add_temp_147; // sfix37_En34
  wire signed [35:0] sum149; // sfix36_En34
  wire signed [35:0] add_signext_296; // sfix36_En34
  wire signed [35:0] add_signext_297; // sfix36_En34
  wire signed [36:0] add_temp_148; // sfix37_En34
  wire signed [35:0] sum150; // sfix36_En34
  wire signed [35:0] add_signext_298; // sfix36_En34
  wire signed [35:0] add_signext_299; // sfix36_En34
  wire signed [36:0] add_temp_149; // sfix37_En34
  wire signed [35:0] sum151; // sfix36_En34
  wire signed [35:0] add_signext_300; // sfix36_En34
  wire signed [35:0] add_signext_301; // sfix36_En34
  wire signed [36:0] add_temp_150; // sfix37_En34
  wire signed [35:0] sum152; // sfix36_En34
  wire signed [35:0] add_signext_302; // sfix36_En34
  wire signed [35:0] add_signext_303; // sfix36_En34
  wire signed [36:0] add_temp_151; // sfix37_En34
  wire signed [35:0] sum153; // sfix36_En34
  wire signed [35:0] add_signext_304; // sfix36_En34
  wire signed [35:0] add_signext_305; // sfix36_En34
  wire signed [36:0] add_temp_152; // sfix37_En34
  wire signed [35:0] sum154; // sfix36_En34
  wire signed [35:0] add_signext_306; // sfix36_En34
  wire signed [35:0] add_signext_307; // sfix36_En34
  wire signed [36:0] add_temp_153; // sfix37_En34
  wire signed [35:0] sum155; // sfix36_En34
  wire signed [35:0] add_signext_308; // sfix36_En34
  wire signed [35:0] add_signext_309; // sfix36_En34
  wire signed [36:0] add_temp_154; // sfix37_En34
  wire signed [35:0] sum156; // sfix36_En34
  wire signed [35:0] add_signext_310; // sfix36_En34
  wire signed [35:0] add_signext_311; // sfix36_En34
  wire signed [36:0] add_temp_155; // sfix37_En34
  wire signed [35:0] sum157; // sfix36_En34
  wire signed [35:0] add_signext_312; // sfix36_En34
  wire signed [35:0] add_signext_313; // sfix36_En34
  wire signed [36:0] add_temp_156; // sfix37_En34
  wire signed [35:0] sum158; // sfix36_En34
  wire signed [35:0] add_signext_314; // sfix36_En34
  wire signed [35:0] add_signext_315; // sfix36_En34
  wire signed [36:0] add_temp_157; // sfix37_En34
  wire signed [35:0] sum159; // sfix36_En34
  wire signed [35:0] add_signext_316; // sfix36_En34
  wire signed [35:0] add_signext_317; // sfix36_En34
  wire signed [36:0] add_temp_158; // sfix37_En34
  wire signed [35:0] sum160; // sfix36_En34
  wire signed [35:0] add_signext_318; // sfix36_En34
  wire signed [35:0] add_signext_319; // sfix36_En34
  wire signed [36:0] add_temp_159; // sfix37_En34
  wire signed [35:0] sum161; // sfix36_En34
  wire signed [35:0] add_signext_320; // sfix36_En34
  wire signed [35:0] add_signext_321; // sfix36_En34
  wire signed [36:0] add_temp_160; // sfix37_En34
  wire signed [35:0] sum162; // sfix36_En34
  wire signed [35:0] add_signext_322; // sfix36_En34
  wire signed [35:0] add_signext_323; // sfix36_En34
  wire signed [36:0] add_temp_161; // sfix37_En34
  wire signed [35:0] sum163; // sfix36_En34
  wire signed [35:0] add_signext_324; // sfix36_En34
  wire signed [35:0] add_signext_325; // sfix36_En34
  wire signed [36:0] add_temp_162; // sfix37_En34
  wire signed [35:0] sum164; // sfix36_En34
  wire signed [35:0] add_signext_326; // sfix36_En34
  wire signed [35:0] add_signext_327; // sfix36_En34
  wire signed [36:0] add_temp_163; // sfix37_En34
  wire signed [35:0] sum165; // sfix36_En34
  wire signed [35:0] add_signext_328; // sfix36_En34
  wire signed [35:0] add_signext_329; // sfix36_En34
  wire signed [36:0] add_temp_164; // sfix37_En34
  wire signed [35:0] sum166; // sfix36_En34
  wire signed [35:0] add_signext_330; // sfix36_En34
  wire signed [35:0] add_signext_331; // sfix36_En34
  wire signed [36:0] add_temp_165; // sfix37_En34
  wire signed [35:0] sum167; // sfix36_En34
  wire signed [35:0] add_signext_332; // sfix36_En34
  wire signed [35:0] add_signext_333; // sfix36_En34
  wire signed [36:0] add_temp_166; // sfix37_En34
  wire signed [35:0] sum168; // sfix36_En34
  wire signed [35:0] add_signext_334; // sfix36_En34
  wire signed [35:0] add_signext_335; // sfix36_En34
  wire signed [36:0] add_temp_167; // sfix37_En34
  wire signed [35:0] sum169; // sfix36_En34
  wire signed [35:0] add_signext_336; // sfix36_En34
  wire signed [35:0] add_signext_337; // sfix36_En34
  wire signed [36:0] add_temp_168; // sfix37_En34
  wire signed [35:0] sum170; // sfix36_En34
  wire signed [35:0] add_signext_338; // sfix36_En34
  wire signed [35:0] add_signext_339; // sfix36_En34
  wire signed [36:0] add_temp_169; // sfix37_En34
  wire signed [35:0] sum171; // sfix36_En34
  wire signed [35:0] add_signext_340; // sfix36_En34
  wire signed [35:0] add_signext_341; // sfix36_En34
  wire signed [36:0] add_temp_170; // sfix37_En34
  wire signed [35:0] sum172; // sfix36_En34
  wire signed [35:0] add_signext_342; // sfix36_En34
  wire signed [35:0] add_signext_343; // sfix36_En34
  wire signed [36:0] add_temp_171; // sfix37_En34
  wire signed [35:0] sum173; // sfix36_En34
  wire signed [35:0] add_signext_344; // sfix36_En34
  wire signed [35:0] add_signext_345; // sfix36_En34
  wire signed [36:0] add_temp_172; // sfix37_En34
  wire signed [35:0] sum174; // sfix36_En34
  wire signed [35:0] add_signext_346; // sfix36_En34
  wire signed [35:0] add_signext_347; // sfix36_En34
  wire signed [36:0] add_temp_173; // sfix37_En34
  wire signed [35:0] sum175; // sfix36_En34
  wire signed [35:0] add_signext_348; // sfix36_En34
  wire signed [35:0] add_signext_349; // sfix36_En34
  wire signed [36:0] add_temp_174; // sfix37_En34
  wire signed [35:0] sum176; // sfix36_En34
  wire signed [35:0] add_signext_350; // sfix36_En34
  wire signed [35:0] add_signext_351; // sfix36_En34
  wire signed [36:0] add_temp_175; // sfix37_En34
  wire signed [35:0] sum177; // sfix36_En34
  wire signed [35:0] add_signext_352; // sfix36_En34
  wire signed [35:0] add_signext_353; // sfix36_En34
  wire signed [36:0] add_temp_176; // sfix37_En34
  wire signed [35:0] sum178; // sfix36_En34
  wire signed [35:0] add_signext_354; // sfix36_En34
  wire signed [35:0] add_signext_355; // sfix36_En34
  wire signed [36:0] add_temp_177; // sfix37_En34
  wire signed [35:0] sum179; // sfix36_En34
  wire signed [35:0] add_signext_356; // sfix36_En34
  wire signed [35:0] add_signext_357; // sfix36_En34
  wire signed [36:0] add_temp_178; // sfix37_En34
  wire signed [35:0] sum180; // sfix36_En34
  wire signed [35:0] add_signext_358; // sfix36_En34
  wire signed [35:0] add_signext_359; // sfix36_En34
  wire signed [36:0] add_temp_179; // sfix37_En34
  wire signed [35:0] sum181; // sfix36_En34
  wire signed [35:0] add_signext_360; // sfix36_En34
  wire signed [35:0] add_signext_361; // sfix36_En34
  wire signed [36:0] add_temp_180; // sfix37_En34
  wire signed [35:0] sum182; // sfix36_En34
  wire signed [35:0] add_signext_362; // sfix36_En34
  wire signed [35:0] add_signext_363; // sfix36_En34
  wire signed [36:0] add_temp_181; // sfix37_En34
  wire signed [35:0] sum183; // sfix36_En34
  wire signed [35:0] add_signext_364; // sfix36_En34
  wire signed [35:0] add_signext_365; // sfix36_En34
  wire signed [36:0] add_temp_182; // sfix37_En34
  wire signed [35:0] sum184; // sfix36_En34
  wire signed [35:0] add_signext_366; // sfix36_En34
  wire signed [35:0] add_signext_367; // sfix36_En34
  wire signed [36:0] add_temp_183; // sfix37_En34
  wire signed [35:0] sum185; // sfix36_En34
  wire signed [35:0] add_signext_368; // sfix36_En34
  wire signed [35:0] add_signext_369; // sfix36_En34
  wire signed [36:0] add_temp_184; // sfix37_En34
  wire signed [35:0] sum186; // sfix36_En34
  wire signed [35:0] add_signext_370; // sfix36_En34
  wire signed [35:0] add_signext_371; // sfix36_En34
  wire signed [36:0] add_temp_185; // sfix37_En34
  wire signed [35:0] sum187; // sfix36_En34
  wire signed [35:0] add_signext_372; // sfix36_En34
  wire signed [35:0] add_signext_373; // sfix36_En34
  wire signed [36:0] add_temp_186; // sfix37_En34
  wire signed [35:0] sum188; // sfix36_En34
  wire signed [35:0] add_signext_374; // sfix36_En34
  wire signed [35:0] add_signext_375; // sfix36_En34
  wire signed [36:0] add_temp_187; // sfix37_En34
  wire signed [35:0] sum189; // sfix36_En34
  wire signed [35:0] add_signext_376; // sfix36_En34
  wire signed [35:0] add_signext_377; // sfix36_En34
  wire signed [36:0] add_temp_188; // sfix37_En34
  wire signed [35:0] sum190; // sfix36_En34
  wire signed [35:0] add_signext_378; // sfix36_En34
  wire signed [35:0] add_signext_379; // sfix36_En34
  wire signed [36:0] add_temp_189; // sfix37_En34
  wire signed [35:0] sum191; // sfix36_En34
  wire signed [35:0] add_signext_380; // sfix36_En34
  wire signed [35:0] add_signext_381; // sfix36_En34
  wire signed [36:0] add_temp_190; // sfix37_En34
  wire signed [35:0] sum192; // sfix36_En34
  wire signed [35:0] add_signext_382; // sfix36_En34
  wire signed [35:0] add_signext_383; // sfix36_En34
  wire signed [36:0] add_temp_191; // sfix37_En34
  wire signed [35:0] sum193; // sfix36_En34
  wire signed [35:0] add_signext_384; // sfix36_En34
  wire signed [35:0] add_signext_385; // sfix36_En34
  wire signed [36:0] add_temp_192; // sfix37_En34
  wire signed [35:0] sum194; // sfix36_En34
  wire signed [35:0] add_signext_386; // sfix36_En34
  wire signed [35:0] add_signext_387; // sfix36_En34
  wire signed [36:0] add_temp_193; // sfix37_En34
  wire signed [35:0] sum195; // sfix36_En34
  wire signed [35:0] add_signext_388; // sfix36_En34
  wire signed [35:0] add_signext_389; // sfix36_En34
  wire signed [36:0] add_temp_194; // sfix37_En34
  wire signed [35:0] sum196; // sfix36_En34
  wire signed [35:0] add_signext_390; // sfix36_En34
  wire signed [35:0] add_signext_391; // sfix36_En34
  wire signed [36:0] add_temp_195; // sfix37_En34
  wire signed [35:0] sum197; // sfix36_En34
  wire signed [35:0] add_signext_392; // sfix36_En34
  wire signed [35:0] add_signext_393; // sfix36_En34
  wire signed [36:0] add_temp_196; // sfix37_En34
  wire signed [35:0] sum198; // sfix36_En34
  wire signed [35:0] add_signext_394; // sfix36_En34
  wire signed [35:0] add_signext_395; // sfix36_En34
  wire signed [36:0] add_temp_197; // sfix37_En34
  wire signed [35:0] sum199; // sfix36_En34
  wire signed [35:0] add_signext_396; // sfix36_En34
  wire signed [35:0] add_signext_397; // sfix36_En34
  wire signed [36:0] add_temp_198; // sfix37_En34
  wire signed [35:0] sum200; // sfix36_En34
  wire signed [35:0] add_signext_398; // sfix36_En34
  wire signed [35:0] add_signext_399; // sfix36_En34
  wire signed [36:0] add_temp_199; // sfix37_En34
  wire signed [35:0] sum201; // sfix36_En34
  wire signed [35:0] add_signext_400; // sfix36_En34
  wire signed [35:0] add_signext_401; // sfix36_En34
  wire signed [36:0] add_temp_200; // sfix37_En34
  wire signed [35:0] sum202; // sfix36_En34
  wire signed [35:0] add_signext_402; // sfix36_En34
  wire signed [35:0] add_signext_403; // sfix36_En34
  wire signed [36:0] add_temp_201; // sfix37_En34
  wire signed [35:0] sum203; // sfix36_En34
  wire signed [35:0] add_signext_404; // sfix36_En34
  wire signed [35:0] add_signext_405; // sfix36_En34
  wire signed [36:0] add_temp_202; // sfix37_En34
  wire signed [35:0] sum204; // sfix36_En34
  wire signed [35:0] add_signext_406; // sfix36_En34
  wire signed [35:0] add_signext_407; // sfix36_En34
  wire signed [36:0] add_temp_203; // sfix37_En34
  wire signed [35:0] sum205; // sfix36_En34
  wire signed [35:0] add_signext_408; // sfix36_En34
  wire signed [35:0] add_signext_409; // sfix36_En34
  wire signed [36:0] add_temp_204; // sfix37_En34
  wire signed [35:0] sum206; // sfix36_En34
  wire signed [35:0] add_signext_410; // sfix36_En34
  wire signed [35:0] add_signext_411; // sfix36_En34
  wire signed [36:0] add_temp_205; // sfix37_En34
  wire signed [35:0] sum207; // sfix36_En34
  wire signed [35:0] add_signext_412; // sfix36_En34
  wire signed [35:0] add_signext_413; // sfix36_En34
  wire signed [36:0] add_temp_206; // sfix37_En34
  wire signed [35:0] sum208; // sfix36_En34
  wire signed [35:0] add_signext_414; // sfix36_En34
  wire signed [35:0] add_signext_415; // sfix36_En34
  wire signed [36:0] add_temp_207; // sfix37_En34
  wire signed [35:0] sum209; // sfix36_En34
  wire signed [35:0] add_signext_416; // sfix36_En34
  wire signed [35:0] add_signext_417; // sfix36_En34
  wire signed [36:0] add_temp_208; // sfix37_En34
  wire signed [35:0] sum210; // sfix36_En34
  wire signed [35:0] add_signext_418; // sfix36_En34
  wire signed [35:0] add_signext_419; // sfix36_En34
  wire signed [36:0] add_temp_209; // sfix37_En34
  wire signed [35:0] sum211; // sfix36_En34
  wire signed [35:0] add_signext_420; // sfix36_En34
  wire signed [35:0] add_signext_421; // sfix36_En34
  wire signed [36:0] add_temp_210; // sfix37_En34
  reg  signed [35:0] output_register; // sfix36_En34

  // Block Statements
  always @( posedge clk or posedge reset)
    begin: Delay_Pipeline_process
      if (reset == 1'b1) begin
        delay_pipeline[0] <= 0;
        delay_pipeline[1] <= 0;
        delay_pipeline[2] <= 0;
        delay_pipeline[3] <= 0;
        delay_pipeline[4] <= 0;
        delay_pipeline[5] <= 0;
        delay_pipeline[6] <= 0;
        delay_pipeline[7] <= 0;
        delay_pipeline[8] <= 0;
        delay_pipeline[9] <= 0;
        delay_pipeline[10] <= 0;
        delay_pipeline[11] <= 0;
        delay_pipeline[12] <= 0;
        delay_pipeline[13] <= 0;
        delay_pipeline[14] <= 0;
        delay_pipeline[15] <= 0;
        delay_pipeline[16] <= 0;
        delay_pipeline[17] <= 0;
        delay_pipeline[18] <= 0;
        delay_pipeline[19] <= 0;
        delay_pipeline[20] <= 0;
        delay_pipeline[21] <= 0;
        delay_pipeline[22] <= 0;
        delay_pipeline[23] <= 0;
        delay_pipeline[24] <= 0;
        delay_pipeline[25] <= 0;
        delay_pipeline[26] <= 0;
        delay_pipeline[27] <= 0;
        delay_pipeline[28] <= 0;
        delay_pipeline[29] <= 0;
        delay_pipeline[30] <= 0;
        delay_pipeline[31] <= 0;
        delay_pipeline[32] <= 0;
        delay_pipeline[33] <= 0;
        delay_pipeline[34] <= 0;
        delay_pipeline[35] <= 0;
        delay_pipeline[36] <= 0;
        delay_pipeline[37] <= 0;
        delay_pipeline[38] <= 0;
        delay_pipeline[39] <= 0;
        delay_pipeline[40] <= 0;
        delay_pipeline[41] <= 0;
        delay_pipeline[42] <= 0;
        delay_pipeline[43] <= 0;
        delay_pipeline[44] <= 0;
        delay_pipeline[45] <= 0;
        delay_pipeline[46] <= 0;
        delay_pipeline[47] <= 0;
        delay_pipeline[48] <= 0;
        delay_pipeline[49] <= 0;
        delay_pipeline[50] <= 0;
        delay_pipeline[51] <= 0;
        delay_pipeline[52] <= 0;
        delay_pipeline[53] <= 0;
        delay_pipeline[54] <= 0;
        delay_pipeline[55] <= 0;
        delay_pipeline[56] <= 0;
        delay_pipeline[57] <= 0;
        delay_pipeline[58] <= 0;
        delay_pipeline[59] <= 0;
        delay_pipeline[60] <= 0;
        delay_pipeline[61] <= 0;
        delay_pipeline[62] <= 0;
        delay_pipeline[63] <= 0;
        delay_pipeline[64] <= 0;
        delay_pipeline[65] <= 0;
        delay_pipeline[66] <= 0;
        delay_pipeline[67] <= 0;
        delay_pipeline[68] <= 0;
        delay_pipeline[69] <= 0;
        delay_pipeline[70] <= 0;
        delay_pipeline[71] <= 0;
        delay_pipeline[72] <= 0;
        delay_pipeline[73] <= 0;
        delay_pipeline[74] <= 0;
        delay_pipeline[75] <= 0;
        delay_pipeline[76] <= 0;
        delay_pipeline[77] <= 0;
        delay_pipeline[78] <= 0;
        delay_pipeline[79] <= 0;
        delay_pipeline[80] <= 0;
        delay_pipeline[81] <= 0;
        delay_pipeline[82] <= 0;
        delay_pipeline[83] <= 0;
        delay_pipeline[84] <= 0;
        delay_pipeline[85] <= 0;
        delay_pipeline[86] <= 0;
        delay_pipeline[87] <= 0;
        delay_pipeline[88] <= 0;
        delay_pipeline[89] <= 0;
        delay_pipeline[90] <= 0;
        delay_pipeline[91] <= 0;
        delay_pipeline[92] <= 0;
        delay_pipeline[93] <= 0;
        delay_pipeline[94] <= 0;
        delay_pipeline[95] <= 0;
        delay_pipeline[96] <= 0;
        delay_pipeline[97] <= 0;
        delay_pipeline[98] <= 0;
        delay_pipeline[99] <= 0;
        delay_pipeline[100] <= 0;
        delay_pipeline[101] <= 0;
        delay_pipeline[102] <= 0;
        delay_pipeline[103] <= 0;
        delay_pipeline[104] <= 0;
        delay_pipeline[105] <= 0;
        delay_pipeline[106] <= 0;
        delay_pipeline[107] <= 0;
        delay_pipeline[108] <= 0;
        delay_pipeline[109] <= 0;
        delay_pipeline[110] <= 0;
        delay_pipeline[111] <= 0;
        delay_pipeline[112] <= 0;
        delay_pipeline[113] <= 0;
        delay_pipeline[114] <= 0;
        delay_pipeline[115] <= 0;
        delay_pipeline[116] <= 0;
        delay_pipeline[117] <= 0;
        delay_pipeline[118] <= 0;
        delay_pipeline[119] <= 0;
        delay_pipeline[120] <= 0;
        delay_pipeline[121] <= 0;
        delay_pipeline[122] <= 0;
        delay_pipeline[123] <= 0;
        delay_pipeline[124] <= 0;
        delay_pipeline[125] <= 0;
        delay_pipeline[126] <= 0;
        delay_pipeline[127] <= 0;
        delay_pipeline[128] <= 0;
        delay_pipeline[129] <= 0;
        delay_pipeline[130] <= 0;
        delay_pipeline[131] <= 0;
        delay_pipeline[132] <= 0;
        delay_pipeline[133] <= 0;
        delay_pipeline[134] <= 0;
        delay_pipeline[135] <= 0;
        delay_pipeline[136] <= 0;
        delay_pipeline[137] <= 0;
        delay_pipeline[138] <= 0;
        delay_pipeline[139] <= 0;
        delay_pipeline[140] <= 0;
        delay_pipeline[141] <= 0;
        delay_pipeline[142] <= 0;
        delay_pipeline[143] <= 0;
        delay_pipeline[144] <= 0;
        delay_pipeline[145] <= 0;
        delay_pipeline[146] <= 0;
        delay_pipeline[147] <= 0;
        delay_pipeline[148] <= 0;
        delay_pipeline[149] <= 0;
        delay_pipeline[150] <= 0;
        delay_pipeline[151] <= 0;
        delay_pipeline[152] <= 0;
        delay_pipeline[153] <= 0;
        delay_pipeline[154] <= 0;
        delay_pipeline[155] <= 0;
        delay_pipeline[156] <= 0;
        delay_pipeline[157] <= 0;
        delay_pipeline[158] <= 0;
        delay_pipeline[159] <= 0;
        delay_pipeline[160] <= 0;
        delay_pipeline[161] <= 0;
        delay_pipeline[162] <= 0;
        delay_pipeline[163] <= 0;
        delay_pipeline[164] <= 0;
        delay_pipeline[165] <= 0;
        delay_pipeline[166] <= 0;
        delay_pipeline[167] <= 0;
        delay_pipeline[168] <= 0;
        delay_pipeline[169] <= 0;
        delay_pipeline[170] <= 0;
        delay_pipeline[171] <= 0;
        delay_pipeline[172] <= 0;
        delay_pipeline[173] <= 0;
        delay_pipeline[174] <= 0;
        delay_pipeline[175] <= 0;
        delay_pipeline[176] <= 0;
        delay_pipeline[177] <= 0;
        delay_pipeline[178] <= 0;
        delay_pipeline[179] <= 0;
        delay_pipeline[180] <= 0;
        delay_pipeline[181] <= 0;
        delay_pipeline[182] <= 0;
        delay_pipeline[183] <= 0;
        delay_pipeline[184] <= 0;
        delay_pipeline[185] <= 0;
        delay_pipeline[186] <= 0;
        delay_pipeline[187] <= 0;
        delay_pipeline[188] <= 0;
        delay_pipeline[189] <= 0;
        delay_pipeline[190] <= 0;
        delay_pipeline[191] <= 0;
        delay_pipeline[192] <= 0;
        delay_pipeline[193] <= 0;
        delay_pipeline[194] <= 0;
        delay_pipeline[195] <= 0;
        delay_pipeline[196] <= 0;
        delay_pipeline[197] <= 0;
        delay_pipeline[198] <= 0;
        delay_pipeline[199] <= 0;
        delay_pipeline[200] <= 0;
        delay_pipeline[201] <= 0;
        delay_pipeline[202] <= 0;
        delay_pipeline[203] <= 0;
        delay_pipeline[204] <= 0;
        delay_pipeline[205] <= 0;
        delay_pipeline[206] <= 0;
        delay_pipeline[207] <= 0;
        delay_pipeline[208] <= 0;
        delay_pipeline[209] <= 0;
        delay_pipeline[210] <= 0;
        delay_pipeline[211] <= 0;
      end
      else begin
        if (clk_enable == 1'b1) begin
          delay_pipeline[0] <= filter_in;
          delay_pipeline[1] <= delay_pipeline[0];
          delay_pipeline[2] <= delay_pipeline[1];
          delay_pipeline[3] <= delay_pipeline[2];
          delay_pipeline[4] <= delay_pipeline[3];
          delay_pipeline[5] <= delay_pipeline[4];
          delay_pipeline[6] <= delay_pipeline[5];
          delay_pipeline[7] <= delay_pipeline[6];
          delay_pipeline[8] <= delay_pipeline[7];
          delay_pipeline[9] <= delay_pipeline[8];
          delay_pipeline[10] <= delay_pipeline[9];
          delay_pipeline[11] <= delay_pipeline[10];
          delay_pipeline[12] <= delay_pipeline[11];
          delay_pipeline[13] <= delay_pipeline[12];
          delay_pipeline[14] <= delay_pipeline[13];
          delay_pipeline[15] <= delay_pipeline[14];
          delay_pipeline[16] <= delay_pipeline[15];
          delay_pipeline[17] <= delay_pipeline[16];
          delay_pipeline[18] <= delay_pipeline[17];
          delay_pipeline[19] <= delay_pipeline[18];
          delay_pipeline[20] <= delay_pipeline[19];
          delay_pipeline[21] <= delay_pipeline[20];
          delay_pipeline[22] <= delay_pipeline[21];
          delay_pipeline[23] <= delay_pipeline[22];
          delay_pipeline[24] <= delay_pipeline[23];
          delay_pipeline[25] <= delay_pipeline[24];
          delay_pipeline[26] <= delay_pipeline[25];
          delay_pipeline[27] <= delay_pipeline[26];
          delay_pipeline[28] <= delay_pipeline[27];
          delay_pipeline[29] <= delay_pipeline[28];
          delay_pipeline[30] <= delay_pipeline[29];
          delay_pipeline[31] <= delay_pipeline[30];
          delay_pipeline[32] <= delay_pipeline[31];
          delay_pipeline[33] <= delay_pipeline[32];
          delay_pipeline[34] <= delay_pipeline[33];
          delay_pipeline[35] <= delay_pipeline[34];
          delay_pipeline[36] <= delay_pipeline[35];
          delay_pipeline[37] <= delay_pipeline[36];
          delay_pipeline[38] <= delay_pipeline[37];
          delay_pipeline[39] <= delay_pipeline[38];
          delay_pipeline[40] <= delay_pipeline[39];
          delay_pipeline[41] <= delay_pipeline[40];
          delay_pipeline[42] <= delay_pipeline[41];
          delay_pipeline[43] <= delay_pipeline[42];
          delay_pipeline[44] <= delay_pipeline[43];
          delay_pipeline[45] <= delay_pipeline[44];
          delay_pipeline[46] <= delay_pipeline[45];
          delay_pipeline[47] <= delay_pipeline[46];
          delay_pipeline[48] <= delay_pipeline[47];
          delay_pipeline[49] <= delay_pipeline[48];
          delay_pipeline[50] <= delay_pipeline[49];
          delay_pipeline[51] <= delay_pipeline[50];
          delay_pipeline[52] <= delay_pipeline[51];
          delay_pipeline[53] <= delay_pipeline[52];
          delay_pipeline[54] <= delay_pipeline[53];
          delay_pipeline[55] <= delay_pipeline[54];
          delay_pipeline[56] <= delay_pipeline[55];
          delay_pipeline[57] <= delay_pipeline[56];
          delay_pipeline[58] <= delay_pipeline[57];
          delay_pipeline[59] <= delay_pipeline[58];
          delay_pipeline[60] <= delay_pipeline[59];
          delay_pipeline[61] <= delay_pipeline[60];
          delay_pipeline[62] <= delay_pipeline[61];
          delay_pipeline[63] <= delay_pipeline[62];
          delay_pipeline[64] <= delay_pipeline[63];
          delay_pipeline[65] <= delay_pipeline[64];
          delay_pipeline[66] <= delay_pipeline[65];
          delay_pipeline[67] <= delay_pipeline[66];
          delay_pipeline[68] <= delay_pipeline[67];
          delay_pipeline[69] <= delay_pipeline[68];
          delay_pipeline[70] <= delay_pipeline[69];
          delay_pipeline[71] <= delay_pipeline[70];
          delay_pipeline[72] <= delay_pipeline[71];
          delay_pipeline[73] <= delay_pipeline[72];
          delay_pipeline[74] <= delay_pipeline[73];
          delay_pipeline[75] <= delay_pipeline[74];
          delay_pipeline[76] <= delay_pipeline[75];
          delay_pipeline[77] <= delay_pipeline[76];
          delay_pipeline[78] <= delay_pipeline[77];
          delay_pipeline[79] <= delay_pipeline[78];
          delay_pipeline[80] <= delay_pipeline[79];
          delay_pipeline[81] <= delay_pipeline[80];
          delay_pipeline[82] <= delay_pipeline[81];
          delay_pipeline[83] <= delay_pipeline[82];
          delay_pipeline[84] <= delay_pipeline[83];
          delay_pipeline[85] <= delay_pipeline[84];
          delay_pipeline[86] <= delay_pipeline[85];
          delay_pipeline[87] <= delay_pipeline[86];
          delay_pipeline[88] <= delay_pipeline[87];
          delay_pipeline[89] <= delay_pipeline[88];
          delay_pipeline[90] <= delay_pipeline[89];
          delay_pipeline[91] <= delay_pipeline[90];
          delay_pipeline[92] <= delay_pipeline[91];
          delay_pipeline[93] <= delay_pipeline[92];
          delay_pipeline[94] <= delay_pipeline[93];
          delay_pipeline[95] <= delay_pipeline[94];
          delay_pipeline[96] <= delay_pipeline[95];
          delay_pipeline[97] <= delay_pipeline[96];
          delay_pipeline[98] <= delay_pipeline[97];
          delay_pipeline[99] <= delay_pipeline[98];
          delay_pipeline[100] <= delay_pipeline[99];
          delay_pipeline[101] <= delay_pipeline[100];
          delay_pipeline[102] <= delay_pipeline[101];
          delay_pipeline[103] <= delay_pipeline[102];
          delay_pipeline[104] <= delay_pipeline[103];
          delay_pipeline[105] <= delay_pipeline[104];
          delay_pipeline[106] <= delay_pipeline[105];
          delay_pipeline[107] <= delay_pipeline[106];
          delay_pipeline[108] <= delay_pipeline[107];
          delay_pipeline[109] <= delay_pipeline[108];
          delay_pipeline[110] <= delay_pipeline[109];
          delay_pipeline[111] <= delay_pipeline[110];
          delay_pipeline[112] <= delay_pipeline[111];
          delay_pipeline[113] <= delay_pipeline[112];
          delay_pipeline[114] <= delay_pipeline[113];
          delay_pipeline[115] <= delay_pipeline[114];
          delay_pipeline[116] <= delay_pipeline[115];
          delay_pipeline[117] <= delay_pipeline[116];
          delay_pipeline[118] <= delay_pipeline[117];
          delay_pipeline[119] <= delay_pipeline[118];
          delay_pipeline[120] <= delay_pipeline[119];
          delay_pipeline[121] <= delay_pipeline[120];
          delay_pipeline[122] <= delay_pipeline[121];
          delay_pipeline[123] <= delay_pipeline[122];
          delay_pipeline[124] <= delay_pipeline[123];
          delay_pipeline[125] <= delay_pipeline[124];
          delay_pipeline[126] <= delay_pipeline[125];
          delay_pipeline[127] <= delay_pipeline[126];
          delay_pipeline[128] <= delay_pipeline[127];
          delay_pipeline[129] <= delay_pipeline[128];
          delay_pipeline[130] <= delay_pipeline[129];
          delay_pipeline[131] <= delay_pipeline[130];
          delay_pipeline[132] <= delay_pipeline[131];
          delay_pipeline[133] <= delay_pipeline[132];
          delay_pipeline[134] <= delay_pipeline[133];
          delay_pipeline[135] <= delay_pipeline[134];
          delay_pipeline[136] <= delay_pipeline[135];
          delay_pipeline[137] <= delay_pipeline[136];
          delay_pipeline[138] <= delay_pipeline[137];
          delay_pipeline[139] <= delay_pipeline[138];
          delay_pipeline[140] <= delay_pipeline[139];
          delay_pipeline[141] <= delay_pipeline[140];
          delay_pipeline[142] <= delay_pipeline[141];
          delay_pipeline[143] <= delay_pipeline[142];
          delay_pipeline[144] <= delay_pipeline[143];
          delay_pipeline[145] <= delay_pipeline[144];
          delay_pipeline[146] <= delay_pipeline[145];
          delay_pipeline[147] <= delay_pipeline[146];
          delay_pipeline[148] <= delay_pipeline[147];
          delay_pipeline[149] <= delay_pipeline[148];
          delay_pipeline[150] <= delay_pipeline[149];
          delay_pipeline[151] <= delay_pipeline[150];
          delay_pipeline[152] <= delay_pipeline[151];
          delay_pipeline[153] <= delay_pipeline[152];
          delay_pipeline[154] <= delay_pipeline[153];
          delay_pipeline[155] <= delay_pipeline[154];
          delay_pipeline[156] <= delay_pipeline[155];
          delay_pipeline[157] <= delay_pipeline[156];
          delay_pipeline[158] <= delay_pipeline[157];
          delay_pipeline[159] <= delay_pipeline[158];
          delay_pipeline[160] <= delay_pipeline[159];
          delay_pipeline[161] <= delay_pipeline[160];
          delay_pipeline[162] <= delay_pipeline[161];
          delay_pipeline[163] <= delay_pipeline[162];
          delay_pipeline[164] <= delay_pipeline[163];
          delay_pipeline[165] <= delay_pipeline[164];
          delay_pipeline[166] <= delay_pipeline[165];
          delay_pipeline[167] <= delay_pipeline[166];
          delay_pipeline[168] <= delay_pipeline[167];
          delay_pipeline[169] <= delay_pipeline[168];
          delay_pipeline[170] <= delay_pipeline[169];
          delay_pipeline[171] <= delay_pipeline[170];
          delay_pipeline[172] <= delay_pipeline[171];
          delay_pipeline[173] <= delay_pipeline[172];
          delay_pipeline[174] <= delay_pipeline[173];
          delay_pipeline[175] <= delay_pipeline[174];
          delay_pipeline[176] <= delay_pipeline[175];
          delay_pipeline[177] <= delay_pipeline[176];
          delay_pipeline[178] <= delay_pipeline[177];
          delay_pipeline[179] <= delay_pipeline[178];
          delay_pipeline[180] <= delay_pipeline[179];
          delay_pipeline[181] <= delay_pipeline[180];
          delay_pipeline[182] <= delay_pipeline[181];
          delay_pipeline[183] <= delay_pipeline[182];
          delay_pipeline[184] <= delay_pipeline[183];
          delay_pipeline[185] <= delay_pipeline[184];
          delay_pipeline[186] <= delay_pipeline[185];
          delay_pipeline[187] <= delay_pipeline[186];
          delay_pipeline[188] <= delay_pipeline[187];
          delay_pipeline[189] <= delay_pipeline[188];
          delay_pipeline[190] <= delay_pipeline[189];
          delay_pipeline[191] <= delay_pipeline[190];
          delay_pipeline[192] <= delay_pipeline[191];
          delay_pipeline[193] <= delay_pipeline[192];
          delay_pipeline[194] <= delay_pipeline[193];
          delay_pipeline[195] <= delay_pipeline[194];
          delay_pipeline[196] <= delay_pipeline[195];
          delay_pipeline[197] <= delay_pipeline[196];
          delay_pipeline[198] <= delay_pipeline[197];
          delay_pipeline[199] <= delay_pipeline[198];
          delay_pipeline[200] <= delay_pipeline[199];
          delay_pipeline[201] <= delay_pipeline[200];
          delay_pipeline[202] <= delay_pipeline[201];
          delay_pipeline[203] <= delay_pipeline[202];
          delay_pipeline[204] <= delay_pipeline[203];
          delay_pipeline[205] <= delay_pipeline[204];
          delay_pipeline[206] <= delay_pipeline[205];
          delay_pipeline[207] <= delay_pipeline[206];
          delay_pipeline[208] <= delay_pipeline[207];
          delay_pipeline[209] <= delay_pipeline[208];
          delay_pipeline[210] <= delay_pipeline[209];
          delay_pipeline[211] <= delay_pipeline[210];
        end
      end
    end // Delay_Pipeline_process


  assign mul_temp = delay_pipeline[211] * coeff212;
  assign product212 = mul_temp[30:0];

  assign mul_temp_1 = delay_pipeline[210] * coeff211;
  assign product211 = mul_temp_1[30:0];

  assign mul_temp_2 = delay_pipeline[209] * coeff210;
  assign product210 = mul_temp_2[30:0];

  assign mul_temp_3 = delay_pipeline[208] * coeff209;
  assign product209 = mul_temp_3[30:0];

  assign mul_temp_4 = delay_pipeline[207] * coeff208;
  assign product208 = mul_temp_4[30:0];

  assign mul_temp_5 = delay_pipeline[206] * coeff207;
  assign product207 = mul_temp_5[30:0];

  assign mul_temp_6 = delay_pipeline[205] * coeff206;
  assign product206 = mul_temp_6[30:0];

  assign mul_temp_7 = delay_pipeline[204] * coeff205;
  assign product205 = mul_temp_7[30:0];

  assign mul_temp_8 = delay_pipeline[203] * coeff204;
  assign product204 = mul_temp_8[30:0];

  assign mul_temp_9 = delay_pipeline[202] * coeff203;
  assign product203 = mul_temp_9[30:0];

  assign mul_temp_10 = delay_pipeline[201] * coeff202;
  assign product202 = mul_temp_10[30:0];

  assign mul_temp_11 = delay_pipeline[200] * coeff201;
  assign product201 = mul_temp_11[30:0];

  assign mul_temp_12 = delay_pipeline[199] * coeff200;
  assign product200 = mul_temp_12[30:0];

  assign mul_temp_13 = delay_pipeline[198] * coeff199;
  assign product199 = mul_temp_13[30:0];

  assign mul_temp_14 = delay_pipeline[197] * coeff198;
  assign product198 = mul_temp_14[30:0];

  assign mul_temp_15 = delay_pipeline[196] * coeff197;
  assign product197 = mul_temp_15[30:0];

  assign mul_temp_16 = delay_pipeline[195] * coeff196;
  assign product196 = mul_temp_16[30:0];

  assign mul_temp_17 = delay_pipeline[194] * coeff195;
  assign product195 = mul_temp_17[30:0];

  assign mul_temp_18 = delay_pipeline[193] * coeff194;
  assign product194 = mul_temp_18[30:0];

  assign mul_temp_19 = delay_pipeline[192] * coeff193;
  assign product193 = mul_temp_19[30:0];

  assign mul_temp_20 = delay_pipeline[191] * coeff192;
  assign product192 = mul_temp_20[30:0];

  assign mul_temp_21 = delay_pipeline[190] * coeff191;
  assign product191 = mul_temp_21[30:0];

  assign mul_temp_22 = delay_pipeline[189] * coeff190;
  assign product190 = mul_temp_22[30:0];

  assign mul_temp_23 = delay_pipeline[188] * coeff189;
  assign product189 = mul_temp_23[30:0];

  assign mul_temp_24 = delay_pipeline[187] * coeff188;
  assign product188 = mul_temp_24[30:0];

  assign mul_temp_25 = delay_pipeline[186] * coeff187;
  assign product187 = mul_temp_25[30:0];

  assign mul_temp_26 = delay_pipeline[185] * coeff186;
  assign product186 = mul_temp_26[30:0];

  assign mul_temp_27 = delay_pipeline[184] * coeff185;
  assign product185 = mul_temp_27[30:0];

  assign mul_temp_28 = delay_pipeline[183] * coeff184;
  assign product184 = mul_temp_28[30:0];

  assign mul_temp_29 = delay_pipeline[182] * coeff183;
  assign product183 = mul_temp_29[30:0];

  assign mul_temp_30 = delay_pipeline[181] * coeff182;
  assign product182 = mul_temp_30[30:0];

  assign mul_temp_31 = delay_pipeline[180] * coeff181;
  assign product181 = mul_temp_31[30:0];

  assign mul_temp_32 = delay_pipeline[179] * coeff180;
  assign product180 = mul_temp_32[30:0];

  assign mul_temp_33 = delay_pipeline[178] * coeff179;
  assign product179 = mul_temp_33[30:0];

  assign mul_temp_34 = delay_pipeline[177] * coeff178;
  assign product178 = mul_temp_34[30:0];

  assign mul_temp_35 = delay_pipeline[176] * coeff177;
  assign product177 = mul_temp_35[30:0];

  assign mul_temp_36 = delay_pipeline[175] * coeff176;
  assign product176 = mul_temp_36[30:0];

  assign mul_temp_37 = delay_pipeline[174] * coeff175;
  assign product175 = mul_temp_37[30:0];

  assign mul_temp_38 = delay_pipeline[173] * coeff174;
  assign product174 = mul_temp_38[30:0];

  assign mul_temp_39 = delay_pipeline[172] * coeff173;
  assign product173 = mul_temp_39[30:0];

  assign mul_temp_40 = delay_pipeline[171] * coeff172;
  assign product172 = mul_temp_40[30:0];

  assign mul_temp_41 = delay_pipeline[170] * coeff171;
  assign product171 = mul_temp_41[30:0];

  assign mul_temp_42 = delay_pipeline[169] * coeff170;
  assign product170 = mul_temp_42[30:0];

  assign mul_temp_43 = delay_pipeline[168] * coeff169;
  assign product169 = mul_temp_43[30:0];

  assign mul_temp_44 = delay_pipeline[167] * coeff168;
  assign product168 = mul_temp_44[30:0];

  assign mul_temp_45 = delay_pipeline[166] * coeff167;
  assign product167 = mul_temp_45[30:0];

  assign mul_temp_46 = delay_pipeline[165] * coeff166;
  assign product166 = mul_temp_46[30:0];

  assign mul_temp_47 = delay_pipeline[164] * coeff165;
  assign product165 = mul_temp_47[30:0];

  assign mul_temp_48 = delay_pipeline[163] * coeff164;
  assign product164 = mul_temp_48[30:0];

  assign mul_temp_49 = delay_pipeline[162] * coeff163;
  assign product163 = mul_temp_49[30:0];

  assign mul_temp_50 = delay_pipeline[161] * coeff162;
  assign product162 = mul_temp_50[30:0];

  assign mul_temp_51 = delay_pipeline[160] * coeff161;
  assign product161 = mul_temp_51[30:0];

  assign mul_temp_52 = delay_pipeline[159] * coeff160;
  assign product160 = mul_temp_52[30:0];

  assign mul_temp_53 = delay_pipeline[158] * coeff159;
  assign product159 = mul_temp_53[30:0];

  assign mul_temp_54 = delay_pipeline[157] * coeff158;
  assign product158 = mul_temp_54[30:0];

  assign mul_temp_55 = delay_pipeline[156] * coeff157;
  assign product157 = mul_temp_55[30:0];

  assign mul_temp_56 = delay_pipeline[155] * coeff156;
  assign product156 = mul_temp_56[30:0];

  assign mul_temp_57 = delay_pipeline[154] * coeff155;
  assign product155 = mul_temp_57[30:0];

  assign mul_temp_58 = delay_pipeline[153] * coeff154;
  assign product154 = mul_temp_58[30:0];

  assign mul_temp_59 = delay_pipeline[152] * coeff153;
  assign product153 = mul_temp_59[30:0];

  assign mul_temp_60 = delay_pipeline[151] * coeff152;
  assign product152 = mul_temp_60[30:0];

  assign mul_temp_61 = delay_pipeline[150] * coeff151;
  assign product151 = mul_temp_61[30:0];

  assign mul_temp_62 = delay_pipeline[149] * coeff150;
  assign product150 = mul_temp_62[30:0];

  assign mul_temp_63 = delay_pipeline[148] * coeff149;
  assign product149 = mul_temp_63[30:0];

  assign mul_temp_64 = delay_pipeline[147] * coeff148;
  assign product148 = mul_temp_64[30:0];

  assign mul_temp_65 = delay_pipeline[146] * coeff147;
  assign product147 = mul_temp_65[30:0];

  assign mul_temp_66 = delay_pipeline[145] * coeff146;
  assign product146 = mul_temp_66[30:0];

  assign mul_temp_67 = delay_pipeline[144] * coeff145;
  assign product145 = mul_temp_67[30:0];

  assign mul_temp_68 = delay_pipeline[143] * coeff144;
  assign product144 = mul_temp_68[30:0];

  assign mul_temp_69 = delay_pipeline[142] * coeff143;
  assign product143 = mul_temp_69[30:0];

  assign mul_temp_70 = delay_pipeline[141] * coeff142;
  assign product142 = mul_temp_70[30:0];

  assign mul_temp_71 = delay_pipeline[140] * coeff141;
  assign product141 = mul_temp_71[30:0];

  assign mul_temp_72 = delay_pipeline[139] * coeff140;
  assign product140 = mul_temp_72[30:0];

  assign mul_temp_73 = delay_pipeline[138] * coeff139;
  assign product139 = mul_temp_73[30:0];

  assign mul_temp_74 = delay_pipeline[137] * coeff138;
  assign product138 = mul_temp_74[30:0];

  assign mul_temp_75 = delay_pipeline[136] * coeff137;
  assign product137 = mul_temp_75[30:0];

  assign mul_temp_76 = delay_pipeline[135] * coeff136;
  assign product136 = mul_temp_76[30:0];

  assign mul_temp_77 = delay_pipeline[134] * coeff135;
  assign product135 = mul_temp_77[30:0];

  assign mul_temp_78 = delay_pipeline[133] * coeff134;
  assign product134 = mul_temp_78[30:0];

  assign mul_temp_79 = delay_pipeline[132] * coeff133;
  assign product133 = mul_temp_79[30:0];

  assign mul_temp_80 = delay_pipeline[131] * coeff132;
  assign product132 = mul_temp_80[30:0];

  assign mul_temp_81 = delay_pipeline[130] * coeff131;
  assign product131 = mul_temp_81[30:0];

  assign mul_temp_82 = delay_pipeline[129] * coeff130;
  assign product130 = mul_temp_82[30:0];

  assign mul_temp_83 = delay_pipeline[128] * coeff129;
  assign product129 = mul_temp_83[30:0];

  assign mul_temp_84 = delay_pipeline[127] * coeff128;
  assign product128 = mul_temp_84[30:0];

  assign mul_temp_85 = delay_pipeline[126] * coeff127;
  assign product127 = mul_temp_85[30:0];

  assign mul_temp_86 = delay_pipeline[125] * coeff126;
  assign product126 = mul_temp_86[30:0];

  assign mul_temp_87 = delay_pipeline[124] * coeff125;
  assign product125 = mul_temp_87[30:0];

  assign mul_temp_88 = delay_pipeline[123] * coeff124;
  assign product124 = mul_temp_88[30:0];

  assign mul_temp_89 = delay_pipeline[122] * coeff123;
  assign product123 = mul_temp_89[30:0];

  assign mul_temp_90 = delay_pipeline[121] * coeff122;
  assign product122 = mul_temp_90[30:0];

  assign mul_temp_91 = delay_pipeline[120] * coeff121;
  assign product121 = mul_temp_91[30:0];

  assign mul_temp_92 = delay_pipeline[119] * coeff120;
  assign product120 = mul_temp_92[30:0];

  assign mul_temp_93 = delay_pipeline[118] * coeff119;
  assign product119 = mul_temp_93[30:0];

  assign mul_temp_94 = delay_pipeline[117] * coeff118;
  assign product118 = mul_temp_94[30:0];

  assign mul_temp_95 = delay_pipeline[116] * coeff117;
  assign product117 = mul_temp_95[30:0];

  assign mul_temp_96 = delay_pipeline[115] * coeff116;
  assign product116 = mul_temp_96[30:0];

  assign mul_temp_97 = delay_pipeline[114] * coeff115;
  assign product115 = mul_temp_97[30:0];

  assign mul_temp_98 = delay_pipeline[113] * coeff114;
  assign product114 = mul_temp_98[30:0];

  assign mul_temp_99 = delay_pipeline[112] * coeff113;
  assign product113 = mul_temp_99[30:0];

  assign mul_temp_100 = delay_pipeline[111] * coeff112;
  assign product112 = mul_temp_100[30:0];

  assign mul_temp_101 = delay_pipeline[110] * coeff111;
  assign product111 = mul_temp_101[30:0];

  assign mul_temp_102 = delay_pipeline[109] * coeff110;
  assign product110 = mul_temp_102[30:0];

  assign mul_temp_103 = delay_pipeline[108] * coeff109;
  assign product109 = mul_temp_103[30:0];

  assign mul_temp_104 = delay_pipeline[107] * coeff108;
  assign product108 = mul_temp_104[30:0];

  assign mul_temp_105 = delay_pipeline[106] * coeff107;
  assign product107 = mul_temp_105[30:0];

  assign mul_temp_106 = delay_pipeline[105] * coeff106;
  assign product106 = mul_temp_106[30:0];

  assign mul_temp_107 = delay_pipeline[104] * coeff105;
  assign product105 = mul_temp_107[30:0];

  assign mul_temp_108 = delay_pipeline[103] * coeff104;
  assign product104 = mul_temp_108[30:0];

  assign mul_temp_109 = delay_pipeline[102] * coeff103;
  assign product103 = mul_temp_109[30:0];

  assign mul_temp_110 = delay_pipeline[101] * coeff102;
  assign product102 = mul_temp_110[30:0];

  assign mul_temp_111 = delay_pipeline[100] * coeff101;
  assign product101 = mul_temp_111[30:0];

  assign mul_temp_112 = delay_pipeline[99] * coeff100;
  assign product100 = mul_temp_112[30:0];

  assign mul_temp_113 = delay_pipeline[98] * coeff99;
  assign product99 = mul_temp_113[30:0];

  assign mul_temp_114 = delay_pipeline[97] * coeff98;
  assign product98 = mul_temp_114[30:0];

  assign mul_temp_115 = delay_pipeline[96] * coeff97;
  assign product97 = mul_temp_115[30:0];

  assign mul_temp_116 = delay_pipeline[95] * coeff96;
  assign product96 = mul_temp_116[30:0];

  assign mul_temp_117 = delay_pipeline[94] * coeff95;
  assign product95 = mul_temp_117[30:0];

  assign mul_temp_118 = delay_pipeline[93] * coeff94;
  assign product94 = mul_temp_118[30:0];

  assign mul_temp_119 = delay_pipeline[92] * coeff93;
  assign product93 = mul_temp_119[30:0];

  assign mul_temp_120 = delay_pipeline[91] * coeff92;
  assign product92 = mul_temp_120[30:0];

  assign mul_temp_121 = delay_pipeline[90] * coeff91;
  assign product91 = mul_temp_121[30:0];

  assign mul_temp_122 = delay_pipeline[89] * coeff90;
  assign product90 = mul_temp_122[30:0];

  assign mul_temp_123 = delay_pipeline[88] * coeff89;
  assign product89 = mul_temp_123[30:0];

  assign mul_temp_124 = delay_pipeline[87] * coeff88;
  assign product88 = mul_temp_124[30:0];

  assign mul_temp_125 = delay_pipeline[86] * coeff87;
  assign product87 = mul_temp_125[30:0];

  assign mul_temp_126 = delay_pipeline[85] * coeff86;
  assign product86 = mul_temp_126[30:0];

  assign mul_temp_127 = delay_pipeline[84] * coeff85;
  assign product85 = mul_temp_127[30:0];

  assign mul_temp_128 = delay_pipeline[83] * coeff84;
  assign product84 = mul_temp_128[30:0];

  assign mul_temp_129 = delay_pipeline[82] * coeff83;
  assign product83 = mul_temp_129[30:0];

  assign mul_temp_130 = delay_pipeline[81] * coeff82;
  assign product82 = mul_temp_130[30:0];

  assign mul_temp_131 = delay_pipeline[80] * coeff81;
  assign product81 = mul_temp_131[30:0];

  assign mul_temp_132 = delay_pipeline[79] * coeff80;
  assign product80 = mul_temp_132[30:0];

  assign mul_temp_133 = delay_pipeline[78] * coeff79;
  assign product79 = mul_temp_133[30:0];

  assign mul_temp_134 = delay_pipeline[77] * coeff78;
  assign product78 = mul_temp_134[30:0];

  assign mul_temp_135 = delay_pipeline[76] * coeff77;
  assign product77 = mul_temp_135[30:0];

  assign mul_temp_136 = delay_pipeline[75] * coeff76;
  assign product76 = mul_temp_136[30:0];

  assign mul_temp_137 = delay_pipeline[74] * coeff75;
  assign product75 = mul_temp_137[30:0];

  assign mul_temp_138 = delay_pipeline[73] * coeff74;
  assign product74 = mul_temp_138[30:0];

  assign mul_temp_139 = delay_pipeline[72] * coeff73;
  assign product73 = mul_temp_139[30:0];

  assign mul_temp_140 = delay_pipeline[71] * coeff72;
  assign product72 = mul_temp_140[30:0];

  assign mul_temp_141 = delay_pipeline[70] * coeff71;
  assign product71 = mul_temp_141[30:0];

  assign mul_temp_142 = delay_pipeline[69] * coeff70;
  assign product70 = mul_temp_142[30:0];

  assign mul_temp_143 = delay_pipeline[68] * coeff69;
  assign product69 = mul_temp_143[30:0];

  assign mul_temp_144 = delay_pipeline[67] * coeff68;
  assign product68 = mul_temp_144[30:0];

  assign mul_temp_145 = delay_pipeline[66] * coeff67;
  assign product67 = mul_temp_145[30:0];

  assign mul_temp_146 = delay_pipeline[65] * coeff66;
  assign product66 = mul_temp_146[30:0];

  assign mul_temp_147 = delay_pipeline[64] * coeff65;
  assign product65 = mul_temp_147[30:0];

  assign mul_temp_148 = delay_pipeline[63] * coeff64;
  assign product64 = mul_temp_148[30:0];

  assign mul_temp_149 = delay_pipeline[62] * coeff63;
  assign product63 = mul_temp_149[30:0];

  assign mul_temp_150 = delay_pipeline[61] * coeff62;
  assign product62 = mul_temp_150[30:0];

  assign mul_temp_151 = delay_pipeline[60] * coeff61;
  assign product61 = mul_temp_151[30:0];

  assign mul_temp_152 = delay_pipeline[59] * coeff60;
  assign product60 = mul_temp_152[30:0];

  assign mul_temp_153 = delay_pipeline[58] * coeff59;
  assign product59 = mul_temp_153[30:0];

  assign mul_temp_154 = delay_pipeline[57] * coeff58;
  assign product58 = mul_temp_154[30:0];

  assign mul_temp_155 = delay_pipeline[56] * coeff57;
  assign product57 = mul_temp_155[30:0];

  assign mul_temp_156 = delay_pipeline[55] * coeff56;
  assign product56 = mul_temp_156[30:0];

  assign mul_temp_157 = delay_pipeline[54] * coeff55;
  assign product55 = mul_temp_157[30:0];

  assign mul_temp_158 = delay_pipeline[53] * coeff54;
  assign product54 = mul_temp_158[30:0];

  assign mul_temp_159 = delay_pipeline[52] * coeff53;
  assign product53 = mul_temp_159[30:0];

  assign mul_temp_160 = delay_pipeline[51] * coeff52;
  assign product52 = mul_temp_160[30:0];

  assign mul_temp_161 = delay_pipeline[50] * coeff51;
  assign product51 = mul_temp_161[30:0];

  assign mul_temp_162 = delay_pipeline[49] * coeff50;
  assign product50 = mul_temp_162[30:0];

  assign mul_temp_163 = delay_pipeline[48] * coeff49;
  assign product49 = mul_temp_163[30:0];

  assign mul_temp_164 = delay_pipeline[47] * coeff48;
  assign product48 = mul_temp_164[30:0];

  assign mul_temp_165 = delay_pipeline[46] * coeff47;
  assign product47 = mul_temp_165[30:0];

  assign mul_temp_166 = delay_pipeline[45] * coeff46;
  assign product46 = mul_temp_166[30:0];

  assign mul_temp_167 = delay_pipeline[44] * coeff45;
  assign product45 = mul_temp_167[30:0];

  assign mul_temp_168 = delay_pipeline[43] * coeff44;
  assign product44 = mul_temp_168[30:0];

  assign mul_temp_169 = delay_pipeline[42] * coeff43;
  assign product43 = mul_temp_169[30:0];

  assign mul_temp_170 = delay_pipeline[41] * coeff42;
  assign product42 = mul_temp_170[30:0];

  assign mul_temp_171 = delay_pipeline[40] * coeff41;
  assign product41 = mul_temp_171[30:0];

  assign mul_temp_172 = delay_pipeline[39] * coeff40;
  assign product40 = mul_temp_172[30:0];

  assign mul_temp_173 = delay_pipeline[38] * coeff39;
  assign product39 = mul_temp_173[30:0];

  assign mul_temp_174 = delay_pipeline[37] * coeff38;
  assign product38 = mul_temp_174[30:0];

  assign mul_temp_175 = delay_pipeline[36] * coeff37;
  assign product37 = mul_temp_175[30:0];

  assign mul_temp_176 = delay_pipeline[35] * coeff36;
  assign product36 = mul_temp_176[30:0];

  assign mul_temp_177 = delay_pipeline[34] * coeff35;
  assign product35 = mul_temp_177[30:0];

  assign mul_temp_178 = delay_pipeline[33] * coeff34;
  assign product34 = mul_temp_178[30:0];

  assign mul_temp_179 = delay_pipeline[32] * coeff33;
  assign product33 = mul_temp_179[30:0];

  assign mul_temp_180 = delay_pipeline[31] * coeff32;
  assign product32 = mul_temp_180[30:0];

  assign mul_temp_181 = delay_pipeline[30] * coeff31;
  assign product31 = mul_temp_181[30:0];

  assign mul_temp_182 = delay_pipeline[29] * coeff30;
  assign product30 = mul_temp_182[30:0];

  assign mul_temp_183 = delay_pipeline[28] * coeff29;
  assign product29 = mul_temp_183[30:0];

  assign mul_temp_184 = delay_pipeline[27] * coeff28;
  assign product28 = mul_temp_184[30:0];

  assign mul_temp_185 = delay_pipeline[26] * coeff27;
  assign product27 = mul_temp_185[30:0];

  assign mul_temp_186 = delay_pipeline[25] * coeff26;
  assign product26 = mul_temp_186[30:0];

  assign mul_temp_187 = delay_pipeline[24] * coeff25;
  assign product25 = mul_temp_187[30:0];

  assign mul_temp_188 = delay_pipeline[23] * coeff24;
  assign product24 = mul_temp_188[30:0];

  assign mul_temp_189 = delay_pipeline[22] * coeff23;
  assign product23 = mul_temp_189[30:0];

  assign mul_temp_190 = delay_pipeline[21] * coeff22;
  assign product22 = mul_temp_190[30:0];

  assign mul_temp_191 = delay_pipeline[20] * coeff21;
  assign product21 = mul_temp_191[30:0];

  assign mul_temp_192 = delay_pipeline[19] * coeff20;
  assign product20 = mul_temp_192[30:0];

  assign mul_temp_193 = delay_pipeline[18] * coeff19;
  assign product19 = mul_temp_193[30:0];

  assign mul_temp_194 = delay_pipeline[17] * coeff18;
  assign product18 = mul_temp_194[30:0];

  assign mul_temp_195 = delay_pipeline[16] * coeff17;
  assign product17 = mul_temp_195[30:0];

  assign mul_temp_196 = delay_pipeline[15] * coeff16;
  assign product16 = mul_temp_196[30:0];

  assign mul_temp_197 = delay_pipeline[14] * coeff15;
  assign product15 = mul_temp_197[30:0];

  assign mul_temp_198 = delay_pipeline[13] * coeff14;
  assign product14 = mul_temp_198[30:0];

  assign mul_temp_199 = delay_pipeline[12] * coeff13;
  assign product13 = mul_temp_199[30:0];

  assign mul_temp_200 = delay_pipeline[11] * coeff12;
  assign product12 = mul_temp_200[30:0];

  assign mul_temp_201 = delay_pipeline[10] * coeff11;
  assign product11 = mul_temp_201[30:0];

  assign mul_temp_202 = delay_pipeline[9] * coeff10;
  assign product10 = mul_temp_202[30:0];

  assign mul_temp_203 = delay_pipeline[8] * coeff9;
  assign product9 = mul_temp_203[30:0];

  assign mul_temp_204 = delay_pipeline[7] * coeff8;
  assign product8 = mul_temp_204[30:0];

  assign mul_temp_205 = delay_pipeline[6] * coeff7;
  assign product7 = mul_temp_205[30:0];

  assign mul_temp_206 = delay_pipeline[5] * coeff6;
  assign product6 = mul_temp_206[30:0];

  assign mul_temp_207 = delay_pipeline[4] * coeff5;
  assign product5 = mul_temp_207[30:0];

  assign mul_temp_208 = delay_pipeline[3] * coeff4;
  assign product4 = mul_temp_208[30:0];

  assign mul_temp_209 = delay_pipeline[2] * coeff3;
  assign product3 = mul_temp_209[30:0];

  assign mul_temp_210 = delay_pipeline[1] * coeff2;
  assign product2 = mul_temp_210[30:0];

  assign product1_cast = $signed({{5{product1[30]}}, product1});

  assign mul_temp_211 = delay_pipeline[0] * coeff1;
  assign product1 = mul_temp_211[30:0];

  assign add_signext = product1_cast;
  assign add_signext_1 = $signed({{5{product2[30]}}, product2});
  assign add_temp = add_signext + add_signext_1;
  assign sum1 = add_temp[35:0];

  assign add_signext_2 = sum1;
  assign add_signext_3 = $signed({{5{product3[30]}}, product3});
  assign add_temp_1 = add_signext_2 + add_signext_3;
  assign sum2 = add_temp_1[35:0];

  assign add_signext_4 = sum2;
  assign add_signext_5 = $signed({{5{product4[30]}}, product4});
  assign add_temp_2 = add_signext_4 + add_signext_5;
  assign sum3 = add_temp_2[35:0];

  assign add_signext_6 = sum3;
  assign add_signext_7 = $signed({{5{product5[30]}}, product5});
  assign add_temp_3 = add_signext_6 + add_signext_7;
  assign sum4 = add_temp_3[35:0];

  assign add_signext_8 = sum4;
  assign add_signext_9 = $signed({{5{product6[30]}}, product6});
  assign add_temp_4 = add_signext_8 + add_signext_9;
  assign sum5 = add_temp_4[35:0];

  assign add_signext_10 = sum5;
  assign add_signext_11 = $signed({{5{product7[30]}}, product7});
  assign add_temp_5 = add_signext_10 + add_signext_11;
  assign sum6 = add_temp_5[35:0];

  assign add_signext_12 = sum6;
  assign add_signext_13 = $signed({{5{product8[30]}}, product8});
  assign add_temp_6 = add_signext_12 + add_signext_13;
  assign sum7 = add_temp_6[35:0];

  assign add_signext_14 = sum7;
  assign add_signext_15 = $signed({{5{product9[30]}}, product9});
  assign add_temp_7 = add_signext_14 + add_signext_15;
  assign sum8 = add_temp_7[35:0];

  assign add_signext_16 = sum8;
  assign add_signext_17 = $signed({{5{product10[30]}}, product10});
  assign add_temp_8 = add_signext_16 + add_signext_17;
  assign sum9 = add_temp_8[35:0];

  assign add_signext_18 = sum9;
  assign add_signext_19 = $signed({{5{product11[30]}}, product11});
  assign add_temp_9 = add_signext_18 + add_signext_19;
  assign sum10 = add_temp_9[35:0];

  assign add_signext_20 = sum10;
  assign add_signext_21 = $signed({{5{product12[30]}}, product12});
  assign add_temp_10 = add_signext_20 + add_signext_21;
  assign sum11 = add_temp_10[35:0];

  assign add_signext_22 = sum11;
  assign add_signext_23 = $signed({{5{product13[30]}}, product13});
  assign add_temp_11 = add_signext_22 + add_signext_23;
  assign sum12 = add_temp_11[35:0];

  assign add_signext_24 = sum12;
  assign add_signext_25 = $signed({{5{product14[30]}}, product14});
  assign add_temp_12 = add_signext_24 + add_signext_25;
  assign sum13 = add_temp_12[35:0];

  assign add_signext_26 = sum13;
  assign add_signext_27 = $signed({{5{product15[30]}}, product15});
  assign add_temp_13 = add_signext_26 + add_signext_27;
  assign sum14 = add_temp_13[35:0];

  assign add_signext_28 = sum14;
  assign add_signext_29 = $signed({{5{product16[30]}}, product16});
  assign add_temp_14 = add_signext_28 + add_signext_29;
  assign sum15 = add_temp_14[35:0];

  assign add_signext_30 = sum15;
  assign add_signext_31 = $signed({{5{product17[30]}}, product17});
  assign add_temp_15 = add_signext_30 + add_signext_31;
  assign sum16 = add_temp_15[35:0];

  assign add_signext_32 = sum16;
  assign add_signext_33 = $signed({{5{product18[30]}}, product18});
  assign add_temp_16 = add_signext_32 + add_signext_33;
  assign sum17 = add_temp_16[35:0];

  assign add_signext_34 = sum17;
  assign add_signext_35 = $signed({{5{product19[30]}}, product19});
  assign add_temp_17 = add_signext_34 + add_signext_35;
  assign sum18 = add_temp_17[35:0];

  assign add_signext_36 = sum18;
  assign add_signext_37 = $signed({{5{product20[30]}}, product20});
  assign add_temp_18 = add_signext_36 + add_signext_37;
  assign sum19 = add_temp_18[35:0];

  assign add_signext_38 = sum19;
  assign add_signext_39 = $signed({{5{product21[30]}}, product21});
  assign add_temp_19 = add_signext_38 + add_signext_39;
  assign sum20 = add_temp_19[35:0];

  assign add_signext_40 = sum20;
  assign add_signext_41 = $signed({{5{product22[30]}}, product22});
  assign add_temp_20 = add_signext_40 + add_signext_41;
  assign sum21 = add_temp_20[35:0];

  assign add_signext_42 = sum21;
  assign add_signext_43 = $signed({{5{product23[30]}}, product23});
  assign add_temp_21 = add_signext_42 + add_signext_43;
  assign sum22 = add_temp_21[35:0];

  assign add_signext_44 = sum22;
  assign add_signext_45 = $signed({{5{product24[30]}}, product24});
  assign add_temp_22 = add_signext_44 + add_signext_45;
  assign sum23 = add_temp_22[35:0];

  assign add_signext_46 = sum23;
  assign add_signext_47 = $signed({{5{product25[30]}}, product25});
  assign add_temp_23 = add_signext_46 + add_signext_47;
  assign sum24 = add_temp_23[35:0];

  assign add_signext_48 = sum24;
  assign add_signext_49 = $signed({{5{product26[30]}}, product26});
  assign add_temp_24 = add_signext_48 + add_signext_49;
  assign sum25 = add_temp_24[35:0];

  assign add_signext_50 = sum25;
  assign add_signext_51 = $signed({{5{product27[30]}}, product27});
  assign add_temp_25 = add_signext_50 + add_signext_51;
  assign sum26 = add_temp_25[35:0];

  assign add_signext_52 = sum26;
  assign add_signext_53 = $signed({{5{product28[30]}}, product28});
  assign add_temp_26 = add_signext_52 + add_signext_53;
  assign sum27 = add_temp_26[35:0];

  assign add_signext_54 = sum27;
  assign add_signext_55 = $signed({{5{product29[30]}}, product29});
  assign add_temp_27 = add_signext_54 + add_signext_55;
  assign sum28 = add_temp_27[35:0];

  assign add_signext_56 = sum28;
  assign add_signext_57 = $signed({{5{product30[30]}}, product30});
  assign add_temp_28 = add_signext_56 + add_signext_57;
  assign sum29 = add_temp_28[35:0];

  assign add_signext_58 = sum29;
  assign add_signext_59 = $signed({{5{product31[30]}}, product31});
  assign add_temp_29 = add_signext_58 + add_signext_59;
  assign sum30 = add_temp_29[35:0];

  assign add_signext_60 = sum30;
  assign add_signext_61 = $signed({{5{product32[30]}}, product32});
  assign add_temp_30 = add_signext_60 + add_signext_61;
  assign sum31 = add_temp_30[35:0];

  assign add_signext_62 = sum31;
  assign add_signext_63 = $signed({{5{product33[30]}}, product33});
  assign add_temp_31 = add_signext_62 + add_signext_63;
  assign sum32 = add_temp_31[35:0];

  assign add_signext_64 = sum32;
  assign add_signext_65 = $signed({{5{product34[30]}}, product34});
  assign add_temp_32 = add_signext_64 + add_signext_65;
  assign sum33 = add_temp_32[35:0];

  assign add_signext_66 = sum33;
  assign add_signext_67 = $signed({{5{product35[30]}}, product35});
  assign add_temp_33 = add_signext_66 + add_signext_67;
  assign sum34 = add_temp_33[35:0];

  assign add_signext_68 = sum34;
  assign add_signext_69 = $signed({{5{product36[30]}}, product36});
  assign add_temp_34 = add_signext_68 + add_signext_69;
  assign sum35 = add_temp_34[35:0];

  assign add_signext_70 = sum35;
  assign add_signext_71 = $signed({{5{product37[30]}}, product37});
  assign add_temp_35 = add_signext_70 + add_signext_71;
  assign sum36 = add_temp_35[35:0];

  assign add_signext_72 = sum36;
  assign add_signext_73 = $signed({{5{product38[30]}}, product38});
  assign add_temp_36 = add_signext_72 + add_signext_73;
  assign sum37 = add_temp_36[35:0];

  assign add_signext_74 = sum37;
  assign add_signext_75 = $signed({{5{product39[30]}}, product39});
  assign add_temp_37 = add_signext_74 + add_signext_75;
  assign sum38 = add_temp_37[35:0];

  assign add_signext_76 = sum38;
  assign add_signext_77 = $signed({{5{product40[30]}}, product40});
  assign add_temp_38 = add_signext_76 + add_signext_77;
  assign sum39 = add_temp_38[35:0];

  assign add_signext_78 = sum39;
  assign add_signext_79 = $signed({{5{product41[30]}}, product41});
  assign add_temp_39 = add_signext_78 + add_signext_79;
  assign sum40 = add_temp_39[35:0];

  assign add_signext_80 = sum40;
  assign add_signext_81 = $signed({{5{product42[30]}}, product42});
  assign add_temp_40 = add_signext_80 + add_signext_81;
  assign sum41 = add_temp_40[35:0];

  assign add_signext_82 = sum41;
  assign add_signext_83 = $signed({{5{product43[30]}}, product43});
  assign add_temp_41 = add_signext_82 + add_signext_83;
  assign sum42 = add_temp_41[35:0];

  assign add_signext_84 = sum42;
  assign add_signext_85 = $signed({{5{product44[30]}}, product44});
  assign add_temp_42 = add_signext_84 + add_signext_85;
  assign sum43 = add_temp_42[35:0];

  assign add_signext_86 = sum43;
  assign add_signext_87 = $signed({{5{product45[30]}}, product45});
  assign add_temp_43 = add_signext_86 + add_signext_87;
  assign sum44 = add_temp_43[35:0];

  assign add_signext_88 = sum44;
  assign add_signext_89 = $signed({{5{product46[30]}}, product46});
  assign add_temp_44 = add_signext_88 + add_signext_89;
  assign sum45 = add_temp_44[35:0];

  assign add_signext_90 = sum45;
  assign add_signext_91 = $signed({{5{product47[30]}}, product47});
  assign add_temp_45 = add_signext_90 + add_signext_91;
  assign sum46 = add_temp_45[35:0];

  assign add_signext_92 = sum46;
  assign add_signext_93 = $signed({{5{product48[30]}}, product48});
  assign add_temp_46 = add_signext_92 + add_signext_93;
  assign sum47 = add_temp_46[35:0];

  assign add_signext_94 = sum47;
  assign add_signext_95 = $signed({{5{product49[30]}}, product49});
  assign add_temp_47 = add_signext_94 + add_signext_95;
  assign sum48 = add_temp_47[35:0];

  assign add_signext_96 = sum48;
  assign add_signext_97 = $signed({{5{product50[30]}}, product50});
  assign add_temp_48 = add_signext_96 + add_signext_97;
  assign sum49 = add_temp_48[35:0];

  assign add_signext_98 = sum49;
  assign add_signext_99 = $signed({{5{product51[30]}}, product51});
  assign add_temp_49 = add_signext_98 + add_signext_99;
  assign sum50 = add_temp_49[35:0];

  assign add_signext_100 = sum50;
  assign add_signext_101 = $signed({{5{product52[30]}}, product52});
  assign add_temp_50 = add_signext_100 + add_signext_101;
  assign sum51 = add_temp_50[35:0];

  assign add_signext_102 = sum51;
  assign add_signext_103 = $signed({{5{product53[30]}}, product53});
  assign add_temp_51 = add_signext_102 + add_signext_103;
  assign sum52 = add_temp_51[35:0];

  assign add_signext_104 = sum52;
  assign add_signext_105 = $signed({{5{product54[30]}}, product54});
  assign add_temp_52 = add_signext_104 + add_signext_105;
  assign sum53 = add_temp_52[35:0];

  assign add_signext_106 = sum53;
  assign add_signext_107 = $signed({{5{product55[30]}}, product55});
  assign add_temp_53 = add_signext_106 + add_signext_107;
  assign sum54 = add_temp_53[35:0];

  assign add_signext_108 = sum54;
  assign add_signext_109 = $signed({{5{product56[30]}}, product56});
  assign add_temp_54 = add_signext_108 + add_signext_109;
  assign sum55 = add_temp_54[35:0];

  assign add_signext_110 = sum55;
  assign add_signext_111 = $signed({{5{product57[30]}}, product57});
  assign add_temp_55 = add_signext_110 + add_signext_111;
  assign sum56 = add_temp_55[35:0];

  assign add_signext_112 = sum56;
  assign add_signext_113 = $signed({{5{product58[30]}}, product58});
  assign add_temp_56 = add_signext_112 + add_signext_113;
  assign sum57 = add_temp_56[35:0];

  assign add_signext_114 = sum57;
  assign add_signext_115 = $signed({{5{product59[30]}}, product59});
  assign add_temp_57 = add_signext_114 + add_signext_115;
  assign sum58 = add_temp_57[35:0];

  assign add_signext_116 = sum58;
  assign add_signext_117 = $signed({{5{product60[30]}}, product60});
  assign add_temp_58 = add_signext_116 + add_signext_117;
  assign sum59 = add_temp_58[35:0];

  assign add_signext_118 = sum59;
  assign add_signext_119 = $signed({{5{product61[30]}}, product61});
  assign add_temp_59 = add_signext_118 + add_signext_119;
  assign sum60 = add_temp_59[35:0];

  assign add_signext_120 = sum60;
  assign add_signext_121 = $signed({{5{product62[30]}}, product62});
  assign add_temp_60 = add_signext_120 + add_signext_121;
  assign sum61 = add_temp_60[35:0];

  assign add_signext_122 = sum61;
  assign add_signext_123 = $signed({{5{product63[30]}}, product63});
  assign add_temp_61 = add_signext_122 + add_signext_123;
  assign sum62 = add_temp_61[35:0];

  assign add_signext_124 = sum62;
  assign add_signext_125 = $signed({{5{product64[30]}}, product64});
  assign add_temp_62 = add_signext_124 + add_signext_125;
  assign sum63 = add_temp_62[35:0];

  assign add_signext_126 = sum63;
  assign add_signext_127 = $signed({{5{product65[30]}}, product65});
  assign add_temp_63 = add_signext_126 + add_signext_127;
  assign sum64 = add_temp_63[35:0];

  assign add_signext_128 = sum64;
  assign add_signext_129 = $signed({{5{product66[30]}}, product66});
  assign add_temp_64 = add_signext_128 + add_signext_129;
  assign sum65 = add_temp_64[35:0];

  assign add_signext_130 = sum65;
  assign add_signext_131 = $signed({{5{product67[30]}}, product67});
  assign add_temp_65 = add_signext_130 + add_signext_131;
  assign sum66 = add_temp_65[35:0];

  assign add_signext_132 = sum66;
  assign add_signext_133 = $signed({{5{product68[30]}}, product68});
  assign add_temp_66 = add_signext_132 + add_signext_133;
  assign sum67 = add_temp_66[35:0];

  assign add_signext_134 = sum67;
  assign add_signext_135 = $signed({{5{product69[30]}}, product69});
  assign add_temp_67 = add_signext_134 + add_signext_135;
  assign sum68 = add_temp_67[35:0];

  assign add_signext_136 = sum68;
  assign add_signext_137 = $signed({{5{product70[30]}}, product70});
  assign add_temp_68 = add_signext_136 + add_signext_137;
  assign sum69 = add_temp_68[35:0];

  assign add_signext_138 = sum69;
  assign add_signext_139 = $signed({{5{product71[30]}}, product71});
  assign add_temp_69 = add_signext_138 + add_signext_139;
  assign sum70 = add_temp_69[35:0];

  assign add_signext_140 = sum70;
  assign add_signext_141 = $signed({{5{product72[30]}}, product72});
  assign add_temp_70 = add_signext_140 + add_signext_141;
  assign sum71 = add_temp_70[35:0];

  assign add_signext_142 = sum71;
  assign add_signext_143 = $signed({{5{product73[30]}}, product73});
  assign add_temp_71 = add_signext_142 + add_signext_143;
  assign sum72 = add_temp_71[35:0];

  assign add_signext_144 = sum72;
  assign add_signext_145 = $signed({{5{product74[30]}}, product74});
  assign add_temp_72 = add_signext_144 + add_signext_145;
  assign sum73 = add_temp_72[35:0];

  assign add_signext_146 = sum73;
  assign add_signext_147 = $signed({{5{product75[30]}}, product75});
  assign add_temp_73 = add_signext_146 + add_signext_147;
  assign sum74 = add_temp_73[35:0];

  assign add_signext_148 = sum74;
  assign add_signext_149 = $signed({{5{product76[30]}}, product76});
  assign add_temp_74 = add_signext_148 + add_signext_149;
  assign sum75 = add_temp_74[35:0];

  assign add_signext_150 = sum75;
  assign add_signext_151 = $signed({{5{product77[30]}}, product77});
  assign add_temp_75 = add_signext_150 + add_signext_151;
  assign sum76 = add_temp_75[35:0];

  assign add_signext_152 = sum76;
  assign add_signext_153 = $signed({{5{product78[30]}}, product78});
  assign add_temp_76 = add_signext_152 + add_signext_153;
  assign sum77 = add_temp_76[35:0];

  assign add_signext_154 = sum77;
  assign add_signext_155 = $signed({{5{product79[30]}}, product79});
  assign add_temp_77 = add_signext_154 + add_signext_155;
  assign sum78 = add_temp_77[35:0];

  assign add_signext_156 = sum78;
  assign add_signext_157 = $signed({{5{product80[30]}}, product80});
  assign add_temp_78 = add_signext_156 + add_signext_157;
  assign sum79 = add_temp_78[35:0];

  assign add_signext_158 = sum79;
  assign add_signext_159 = $signed({{5{product81[30]}}, product81});
  assign add_temp_79 = add_signext_158 + add_signext_159;
  assign sum80 = add_temp_79[35:0];

  assign add_signext_160 = sum80;
  assign add_signext_161 = $signed({{5{product82[30]}}, product82});
  assign add_temp_80 = add_signext_160 + add_signext_161;
  assign sum81 = add_temp_80[35:0];

  assign add_signext_162 = sum81;
  assign add_signext_163 = $signed({{5{product83[30]}}, product83});
  assign add_temp_81 = add_signext_162 + add_signext_163;
  assign sum82 = add_temp_81[35:0];

  assign add_signext_164 = sum82;
  assign add_signext_165 = $signed({{5{product84[30]}}, product84});
  assign add_temp_82 = add_signext_164 + add_signext_165;
  assign sum83 = add_temp_82[35:0];

  assign add_signext_166 = sum83;
  assign add_signext_167 = $signed({{5{product85[30]}}, product85});
  assign add_temp_83 = add_signext_166 + add_signext_167;
  assign sum84 = add_temp_83[35:0];

  assign add_signext_168 = sum84;
  assign add_signext_169 = $signed({{5{product86[30]}}, product86});
  assign add_temp_84 = add_signext_168 + add_signext_169;
  assign sum85 = add_temp_84[35:0];

  assign add_signext_170 = sum85;
  assign add_signext_171 = $signed({{5{product87[30]}}, product87});
  assign add_temp_85 = add_signext_170 + add_signext_171;
  assign sum86 = add_temp_85[35:0];

  assign add_signext_172 = sum86;
  assign add_signext_173 = $signed({{5{product88[30]}}, product88});
  assign add_temp_86 = add_signext_172 + add_signext_173;
  assign sum87 = add_temp_86[35:0];

  assign add_signext_174 = sum87;
  assign add_signext_175 = $signed({{5{product89[30]}}, product89});
  assign add_temp_87 = add_signext_174 + add_signext_175;
  assign sum88 = add_temp_87[35:0];

  assign add_signext_176 = sum88;
  assign add_signext_177 = $signed({{5{product90[30]}}, product90});
  assign add_temp_88 = add_signext_176 + add_signext_177;
  assign sum89 = add_temp_88[35:0];

  assign add_signext_178 = sum89;
  assign add_signext_179 = $signed({{5{product91[30]}}, product91});
  assign add_temp_89 = add_signext_178 + add_signext_179;
  assign sum90 = add_temp_89[35:0];

  assign add_signext_180 = sum90;
  assign add_signext_181 = $signed({{5{product92[30]}}, product92});
  assign add_temp_90 = add_signext_180 + add_signext_181;
  assign sum91 = add_temp_90[35:0];

  assign add_signext_182 = sum91;
  assign add_signext_183 = $signed({{5{product93[30]}}, product93});
  assign add_temp_91 = add_signext_182 + add_signext_183;
  assign sum92 = add_temp_91[35:0];

  assign add_signext_184 = sum92;
  assign add_signext_185 = $signed({{5{product94[30]}}, product94});
  assign add_temp_92 = add_signext_184 + add_signext_185;
  assign sum93 = add_temp_92[35:0];

  assign add_signext_186 = sum93;
  assign add_signext_187 = $signed({{5{product95[30]}}, product95});
  assign add_temp_93 = add_signext_186 + add_signext_187;
  assign sum94 = add_temp_93[35:0];

  assign add_signext_188 = sum94;
  assign add_signext_189 = $signed({{5{product96[30]}}, product96});
  assign add_temp_94 = add_signext_188 + add_signext_189;
  assign sum95 = add_temp_94[35:0];

  assign add_signext_190 = sum95;
  assign add_signext_191 = $signed({{5{product97[30]}}, product97});
  assign add_temp_95 = add_signext_190 + add_signext_191;
  assign sum96 = add_temp_95[35:0];

  assign add_signext_192 = sum96;
  assign add_signext_193 = $signed({{5{product98[30]}}, product98});
  assign add_temp_96 = add_signext_192 + add_signext_193;
  assign sum97 = add_temp_96[35:0];

  assign add_signext_194 = sum97;
  assign add_signext_195 = $signed({{5{product99[30]}}, product99});
  assign add_temp_97 = add_signext_194 + add_signext_195;
  assign sum98 = add_temp_97[35:0];

  assign add_signext_196 = sum98;
  assign add_signext_197 = $signed({{5{product100[30]}}, product100});
  assign add_temp_98 = add_signext_196 + add_signext_197;
  assign sum99 = add_temp_98[35:0];

  assign add_signext_198 = sum99;
  assign add_signext_199 = $signed({{5{product101[30]}}, product101});
  assign add_temp_99 = add_signext_198 + add_signext_199;
  assign sum100 = add_temp_99[35:0];

  assign add_signext_200 = sum100;
  assign add_signext_201 = $signed({{5{product102[30]}}, product102});
  assign add_temp_100 = add_signext_200 + add_signext_201;
  assign sum101 = add_temp_100[35:0];

  assign add_signext_202 = sum101;
  assign add_signext_203 = $signed({{5{product103[30]}}, product103});
  assign add_temp_101 = add_signext_202 + add_signext_203;
  assign sum102 = add_temp_101[35:0];

  assign add_signext_204 = sum102;
  assign add_signext_205 = $signed({{5{product104[30]}}, product104});
  assign add_temp_102 = add_signext_204 + add_signext_205;
  assign sum103 = add_temp_102[35:0];

  assign add_signext_206 = sum103;
  assign add_signext_207 = $signed({{5{product105[30]}}, product105});
  assign add_temp_103 = add_signext_206 + add_signext_207;
  assign sum104 = add_temp_103[35:0];

  assign add_signext_208 = sum104;
  assign add_signext_209 = $signed({{5{product106[30]}}, product106});
  assign add_temp_104 = add_signext_208 + add_signext_209;
  assign sum105 = add_temp_104[35:0];

  assign add_signext_210 = sum105;
  assign add_signext_211 = $signed({{5{product107[30]}}, product107});
  assign add_temp_105 = add_signext_210 + add_signext_211;
  assign sum106 = add_temp_105[35:0];

  assign add_signext_212 = sum106;
  assign add_signext_213 = $signed({{5{product108[30]}}, product108});
  assign add_temp_106 = add_signext_212 + add_signext_213;
  assign sum107 = add_temp_106[35:0];

  assign add_signext_214 = sum107;
  assign add_signext_215 = $signed({{5{product109[30]}}, product109});
  assign add_temp_107 = add_signext_214 + add_signext_215;
  assign sum108 = add_temp_107[35:0];

  assign add_signext_216 = sum108;
  assign add_signext_217 = $signed({{5{product110[30]}}, product110});
  assign add_temp_108 = add_signext_216 + add_signext_217;
  assign sum109 = add_temp_108[35:0];

  assign add_signext_218 = sum109;
  assign add_signext_219 = $signed({{5{product111[30]}}, product111});
  assign add_temp_109 = add_signext_218 + add_signext_219;
  assign sum110 = add_temp_109[35:0];

  assign add_signext_220 = sum110;
  assign add_signext_221 = $signed({{5{product112[30]}}, product112});
  assign add_temp_110 = add_signext_220 + add_signext_221;
  assign sum111 = add_temp_110[35:0];

  assign add_signext_222 = sum111;
  assign add_signext_223 = $signed({{5{product113[30]}}, product113});
  assign add_temp_111 = add_signext_222 + add_signext_223;
  assign sum112 = add_temp_111[35:0];

  assign add_signext_224 = sum112;
  assign add_signext_225 = $signed({{5{product114[30]}}, product114});
  assign add_temp_112 = add_signext_224 + add_signext_225;
  assign sum113 = add_temp_112[35:0];

  assign add_signext_226 = sum113;
  assign add_signext_227 = $signed({{5{product115[30]}}, product115});
  assign add_temp_113 = add_signext_226 + add_signext_227;
  assign sum114 = add_temp_113[35:0];

  assign add_signext_228 = sum114;
  assign add_signext_229 = $signed({{5{product116[30]}}, product116});
  assign add_temp_114 = add_signext_228 + add_signext_229;
  assign sum115 = add_temp_114[35:0];

  assign add_signext_230 = sum115;
  assign add_signext_231 = $signed({{5{product117[30]}}, product117});
  assign add_temp_115 = add_signext_230 + add_signext_231;
  assign sum116 = add_temp_115[35:0];

  assign add_signext_232 = sum116;
  assign add_signext_233 = $signed({{5{product118[30]}}, product118});
  assign add_temp_116 = add_signext_232 + add_signext_233;
  assign sum117 = add_temp_116[35:0];

  assign add_signext_234 = sum117;
  assign add_signext_235 = $signed({{5{product119[30]}}, product119});
  assign add_temp_117 = add_signext_234 + add_signext_235;
  assign sum118 = add_temp_117[35:0];

  assign add_signext_236 = sum118;
  assign add_signext_237 = $signed({{5{product120[30]}}, product120});
  assign add_temp_118 = add_signext_236 + add_signext_237;
  assign sum119 = add_temp_118[35:0];

  assign add_signext_238 = sum119;
  assign add_signext_239 = $signed({{5{product121[30]}}, product121});
  assign add_temp_119 = add_signext_238 + add_signext_239;
  assign sum120 = add_temp_119[35:0];

  assign add_signext_240 = sum120;
  assign add_signext_241 = $signed({{5{product122[30]}}, product122});
  assign add_temp_120 = add_signext_240 + add_signext_241;
  assign sum121 = add_temp_120[35:0];

  assign add_signext_242 = sum121;
  assign add_signext_243 = $signed({{5{product123[30]}}, product123});
  assign add_temp_121 = add_signext_242 + add_signext_243;
  assign sum122 = add_temp_121[35:0];

  assign add_signext_244 = sum122;
  assign add_signext_245 = $signed({{5{product124[30]}}, product124});
  assign add_temp_122 = add_signext_244 + add_signext_245;
  assign sum123 = add_temp_122[35:0];

  assign add_signext_246 = sum123;
  assign add_signext_247 = $signed({{5{product125[30]}}, product125});
  assign add_temp_123 = add_signext_246 + add_signext_247;
  assign sum124 = add_temp_123[35:0];

  assign add_signext_248 = sum124;
  assign add_signext_249 = $signed({{5{product126[30]}}, product126});
  assign add_temp_124 = add_signext_248 + add_signext_249;
  assign sum125 = add_temp_124[35:0];

  assign add_signext_250 = sum125;
  assign add_signext_251 = $signed({{5{product127[30]}}, product127});
  assign add_temp_125 = add_signext_250 + add_signext_251;
  assign sum126 = add_temp_125[35:0];

  assign add_signext_252 = sum126;
  assign add_signext_253 = $signed({{5{product128[30]}}, product128});
  assign add_temp_126 = add_signext_252 + add_signext_253;
  assign sum127 = add_temp_126[35:0];

  assign add_signext_254 = sum127;
  assign add_signext_255 = $signed({{5{product129[30]}}, product129});
  assign add_temp_127 = add_signext_254 + add_signext_255;
  assign sum128 = add_temp_127[35:0];

  assign add_signext_256 = sum128;
  assign add_signext_257 = $signed({{5{product130[30]}}, product130});
  assign add_temp_128 = add_signext_256 + add_signext_257;
  assign sum129 = add_temp_128[35:0];

  assign add_signext_258 = sum129;
  assign add_signext_259 = $signed({{5{product131[30]}}, product131});
  assign add_temp_129 = add_signext_258 + add_signext_259;
  assign sum130 = add_temp_129[35:0];

  assign add_signext_260 = sum130;
  assign add_signext_261 = $signed({{5{product132[30]}}, product132});
  assign add_temp_130 = add_signext_260 + add_signext_261;
  assign sum131 = add_temp_130[35:0];

  assign add_signext_262 = sum131;
  assign add_signext_263 = $signed({{5{product133[30]}}, product133});
  assign add_temp_131 = add_signext_262 + add_signext_263;
  assign sum132 = add_temp_131[35:0];

  assign add_signext_264 = sum132;
  assign add_signext_265 = $signed({{5{product134[30]}}, product134});
  assign add_temp_132 = add_signext_264 + add_signext_265;
  assign sum133 = add_temp_132[35:0];

  assign add_signext_266 = sum133;
  assign add_signext_267 = $signed({{5{product135[30]}}, product135});
  assign add_temp_133 = add_signext_266 + add_signext_267;
  assign sum134 = add_temp_133[35:0];

  assign add_signext_268 = sum134;
  assign add_signext_269 = $signed({{5{product136[30]}}, product136});
  assign add_temp_134 = add_signext_268 + add_signext_269;
  assign sum135 = add_temp_134[35:0];

  assign add_signext_270 = sum135;
  assign add_signext_271 = $signed({{5{product137[30]}}, product137});
  assign add_temp_135 = add_signext_270 + add_signext_271;
  assign sum136 = add_temp_135[35:0];

  assign add_signext_272 = sum136;
  assign add_signext_273 = $signed({{5{product138[30]}}, product138});
  assign add_temp_136 = add_signext_272 + add_signext_273;
  assign sum137 = add_temp_136[35:0];

  assign add_signext_274 = sum137;
  assign add_signext_275 = $signed({{5{product139[30]}}, product139});
  assign add_temp_137 = add_signext_274 + add_signext_275;
  assign sum138 = add_temp_137[35:0];

  assign add_signext_276 = sum138;
  assign add_signext_277 = $signed({{5{product140[30]}}, product140});
  assign add_temp_138 = add_signext_276 + add_signext_277;
  assign sum139 = add_temp_138[35:0];

  assign add_signext_278 = sum139;
  assign add_signext_279 = $signed({{5{product141[30]}}, product141});
  assign add_temp_139 = add_signext_278 + add_signext_279;
  assign sum140 = add_temp_139[35:0];

  assign add_signext_280 = sum140;
  assign add_signext_281 = $signed({{5{product142[30]}}, product142});
  assign add_temp_140 = add_signext_280 + add_signext_281;
  assign sum141 = add_temp_140[35:0];

  assign add_signext_282 = sum141;
  assign add_signext_283 = $signed({{5{product143[30]}}, product143});
  assign add_temp_141 = add_signext_282 + add_signext_283;
  assign sum142 = add_temp_141[35:0];

  assign add_signext_284 = sum142;
  assign add_signext_285 = $signed({{5{product144[30]}}, product144});
  assign add_temp_142 = add_signext_284 + add_signext_285;
  assign sum143 = add_temp_142[35:0];

  assign add_signext_286 = sum143;
  assign add_signext_287 = $signed({{5{product145[30]}}, product145});
  assign add_temp_143 = add_signext_286 + add_signext_287;
  assign sum144 = add_temp_143[35:0];

  assign add_signext_288 = sum144;
  assign add_signext_289 = $signed({{5{product146[30]}}, product146});
  assign add_temp_144 = add_signext_288 + add_signext_289;
  assign sum145 = add_temp_144[35:0];

  assign add_signext_290 = sum145;
  assign add_signext_291 = $signed({{5{product147[30]}}, product147});
  assign add_temp_145 = add_signext_290 + add_signext_291;
  assign sum146 = add_temp_145[35:0];

  assign add_signext_292 = sum146;
  assign add_signext_293 = $signed({{5{product148[30]}}, product148});
  assign add_temp_146 = add_signext_292 + add_signext_293;
  assign sum147 = add_temp_146[35:0];

  assign add_signext_294 = sum147;
  assign add_signext_295 = $signed({{5{product149[30]}}, product149});
  assign add_temp_147 = add_signext_294 + add_signext_295;
  assign sum148 = add_temp_147[35:0];

  assign add_signext_296 = sum148;
  assign add_signext_297 = $signed({{5{product150[30]}}, product150});
  assign add_temp_148 = add_signext_296 + add_signext_297;
  assign sum149 = add_temp_148[35:0];

  assign add_signext_298 = sum149;
  assign add_signext_299 = $signed({{5{product151[30]}}, product151});
  assign add_temp_149 = add_signext_298 + add_signext_299;
  assign sum150 = add_temp_149[35:0];

  assign add_signext_300 = sum150;
  assign add_signext_301 = $signed({{5{product152[30]}}, product152});
  assign add_temp_150 = add_signext_300 + add_signext_301;
  assign sum151 = add_temp_150[35:0];

  assign add_signext_302 = sum151;
  assign add_signext_303 = $signed({{5{product153[30]}}, product153});
  assign add_temp_151 = add_signext_302 + add_signext_303;
  assign sum152 = add_temp_151[35:0];

  assign add_signext_304 = sum152;
  assign add_signext_305 = $signed({{5{product154[30]}}, product154});
  assign add_temp_152 = add_signext_304 + add_signext_305;
  assign sum153 = add_temp_152[35:0];

  assign add_signext_306 = sum153;
  assign add_signext_307 = $signed({{5{product155[30]}}, product155});
  assign add_temp_153 = add_signext_306 + add_signext_307;
  assign sum154 = add_temp_153[35:0];

  assign add_signext_308 = sum154;
  assign add_signext_309 = $signed({{5{product156[30]}}, product156});
  assign add_temp_154 = add_signext_308 + add_signext_309;
  assign sum155 = add_temp_154[35:0];

  assign add_signext_310 = sum155;
  assign add_signext_311 = $signed({{5{product157[30]}}, product157});
  assign add_temp_155 = add_signext_310 + add_signext_311;
  assign sum156 = add_temp_155[35:0];

  assign add_signext_312 = sum156;
  assign add_signext_313 = $signed({{5{product158[30]}}, product158});
  assign add_temp_156 = add_signext_312 + add_signext_313;
  assign sum157 = add_temp_156[35:0];

  assign add_signext_314 = sum157;
  assign add_signext_315 = $signed({{5{product159[30]}}, product159});
  assign add_temp_157 = add_signext_314 + add_signext_315;
  assign sum158 = add_temp_157[35:0];

  assign add_signext_316 = sum158;
  assign add_signext_317 = $signed({{5{product160[30]}}, product160});
  assign add_temp_158 = add_signext_316 + add_signext_317;
  assign sum159 = add_temp_158[35:0];

  assign add_signext_318 = sum159;
  assign add_signext_319 = $signed({{5{product161[30]}}, product161});
  assign add_temp_159 = add_signext_318 + add_signext_319;
  assign sum160 = add_temp_159[35:0];

  assign add_signext_320 = sum160;
  assign add_signext_321 = $signed({{5{product162[30]}}, product162});
  assign add_temp_160 = add_signext_320 + add_signext_321;
  assign sum161 = add_temp_160[35:0];

  assign add_signext_322 = sum161;
  assign add_signext_323 = $signed({{5{product163[30]}}, product163});
  assign add_temp_161 = add_signext_322 + add_signext_323;
  assign sum162 = add_temp_161[35:0];

  assign add_signext_324 = sum162;
  assign add_signext_325 = $signed({{5{product164[30]}}, product164});
  assign add_temp_162 = add_signext_324 + add_signext_325;
  assign sum163 = add_temp_162[35:0];

  assign add_signext_326 = sum163;
  assign add_signext_327 = $signed({{5{product165[30]}}, product165});
  assign add_temp_163 = add_signext_326 + add_signext_327;
  assign sum164 = add_temp_163[35:0];

  assign add_signext_328 = sum164;
  assign add_signext_329 = $signed({{5{product166[30]}}, product166});
  assign add_temp_164 = add_signext_328 + add_signext_329;
  assign sum165 = add_temp_164[35:0];

  assign add_signext_330 = sum165;
  assign add_signext_331 = $signed({{5{product167[30]}}, product167});
  assign add_temp_165 = add_signext_330 + add_signext_331;
  assign sum166 = add_temp_165[35:0];

  assign add_signext_332 = sum166;
  assign add_signext_333 = $signed({{5{product168[30]}}, product168});
  assign add_temp_166 = add_signext_332 + add_signext_333;
  assign sum167 = add_temp_166[35:0];

  assign add_signext_334 = sum167;
  assign add_signext_335 = $signed({{5{product169[30]}}, product169});
  assign add_temp_167 = add_signext_334 + add_signext_335;
  assign sum168 = add_temp_167[35:0];

  assign add_signext_336 = sum168;
  assign add_signext_337 = $signed({{5{product170[30]}}, product170});
  assign add_temp_168 = add_signext_336 + add_signext_337;
  assign sum169 = add_temp_168[35:0];

  assign add_signext_338 = sum169;
  assign add_signext_339 = $signed({{5{product171[30]}}, product171});
  assign add_temp_169 = add_signext_338 + add_signext_339;
  assign sum170 = add_temp_169[35:0];

  assign add_signext_340 = sum170;
  assign add_signext_341 = $signed({{5{product172[30]}}, product172});
  assign add_temp_170 = add_signext_340 + add_signext_341;
  assign sum171 = add_temp_170[35:0];

  assign add_signext_342 = sum171;
  assign add_signext_343 = $signed({{5{product173[30]}}, product173});
  assign add_temp_171 = add_signext_342 + add_signext_343;
  assign sum172 = add_temp_171[35:0];

  assign add_signext_344 = sum172;
  assign add_signext_345 = $signed({{5{product174[30]}}, product174});
  assign add_temp_172 = add_signext_344 + add_signext_345;
  assign sum173 = add_temp_172[35:0];

  assign add_signext_346 = sum173;
  assign add_signext_347 = $signed({{5{product175[30]}}, product175});
  assign add_temp_173 = add_signext_346 + add_signext_347;
  assign sum174 = add_temp_173[35:0];

  assign add_signext_348 = sum174;
  assign add_signext_349 = $signed({{5{product176[30]}}, product176});
  assign add_temp_174 = add_signext_348 + add_signext_349;
  assign sum175 = add_temp_174[35:0];

  assign add_signext_350 = sum175;
  assign add_signext_351 = $signed({{5{product177[30]}}, product177});
  assign add_temp_175 = add_signext_350 + add_signext_351;
  assign sum176 = add_temp_175[35:0];

  assign add_signext_352 = sum176;
  assign add_signext_353 = $signed({{5{product178[30]}}, product178});
  assign add_temp_176 = add_signext_352 + add_signext_353;
  assign sum177 = add_temp_176[35:0];

  assign add_signext_354 = sum177;
  assign add_signext_355 = $signed({{5{product179[30]}}, product179});
  assign add_temp_177 = add_signext_354 + add_signext_355;
  assign sum178 = add_temp_177[35:0];

  assign add_signext_356 = sum178;
  assign add_signext_357 = $signed({{5{product180[30]}}, product180});
  assign add_temp_178 = add_signext_356 + add_signext_357;
  assign sum179 = add_temp_178[35:0];

  assign add_signext_358 = sum179;
  assign add_signext_359 = $signed({{5{product181[30]}}, product181});
  assign add_temp_179 = add_signext_358 + add_signext_359;
  assign sum180 = add_temp_179[35:0];

  assign add_signext_360 = sum180;
  assign add_signext_361 = $signed({{5{product182[30]}}, product182});
  assign add_temp_180 = add_signext_360 + add_signext_361;
  assign sum181 = add_temp_180[35:0];

  assign add_signext_362 = sum181;
  assign add_signext_363 = $signed({{5{product183[30]}}, product183});
  assign add_temp_181 = add_signext_362 + add_signext_363;
  assign sum182 = add_temp_181[35:0];

  assign add_signext_364 = sum182;
  assign add_signext_365 = $signed({{5{product184[30]}}, product184});
  assign add_temp_182 = add_signext_364 + add_signext_365;
  assign sum183 = add_temp_182[35:0];

  assign add_signext_366 = sum183;
  assign add_signext_367 = $signed({{5{product185[30]}}, product185});
  assign add_temp_183 = add_signext_366 + add_signext_367;
  assign sum184 = add_temp_183[35:0];

  assign add_signext_368 = sum184;
  assign add_signext_369 = $signed({{5{product186[30]}}, product186});
  assign add_temp_184 = add_signext_368 + add_signext_369;
  assign sum185 = add_temp_184[35:0];

  assign add_signext_370 = sum185;
  assign add_signext_371 = $signed({{5{product187[30]}}, product187});
  assign add_temp_185 = add_signext_370 + add_signext_371;
  assign sum186 = add_temp_185[35:0];

  assign add_signext_372 = sum186;
  assign add_signext_373 = $signed({{5{product188[30]}}, product188});
  assign add_temp_186 = add_signext_372 + add_signext_373;
  assign sum187 = add_temp_186[35:0];

  assign add_signext_374 = sum187;
  assign add_signext_375 = $signed({{5{product189[30]}}, product189});
  assign add_temp_187 = add_signext_374 + add_signext_375;
  assign sum188 = add_temp_187[35:0];

  assign add_signext_376 = sum188;
  assign add_signext_377 = $signed({{5{product190[30]}}, product190});
  assign add_temp_188 = add_signext_376 + add_signext_377;
  assign sum189 = add_temp_188[35:0];

  assign add_signext_378 = sum189;
  assign add_signext_379 = $signed({{5{product191[30]}}, product191});
  assign add_temp_189 = add_signext_378 + add_signext_379;
  assign sum190 = add_temp_189[35:0];

  assign add_signext_380 = sum190;
  assign add_signext_381 = $signed({{5{product192[30]}}, product192});
  assign add_temp_190 = add_signext_380 + add_signext_381;
  assign sum191 = add_temp_190[35:0];

  assign add_signext_382 = sum191;
  assign add_signext_383 = $signed({{5{product193[30]}}, product193});
  assign add_temp_191 = add_signext_382 + add_signext_383;
  assign sum192 = add_temp_191[35:0];

  assign add_signext_384 = sum192;
  assign add_signext_385 = $signed({{5{product194[30]}}, product194});
  assign add_temp_192 = add_signext_384 + add_signext_385;
  assign sum193 = add_temp_192[35:0];

  assign add_signext_386 = sum193;
  assign add_signext_387 = $signed({{5{product195[30]}}, product195});
  assign add_temp_193 = add_signext_386 + add_signext_387;
  assign sum194 = add_temp_193[35:0];

  assign add_signext_388 = sum194;
  assign add_signext_389 = $signed({{5{product196[30]}}, product196});
  assign add_temp_194 = add_signext_388 + add_signext_389;
  assign sum195 = add_temp_194[35:0];

  assign add_signext_390 = sum195;
  assign add_signext_391 = $signed({{5{product197[30]}}, product197});
  assign add_temp_195 = add_signext_390 + add_signext_391;
  assign sum196 = add_temp_195[35:0];

  assign add_signext_392 = sum196;
  assign add_signext_393 = $signed({{5{product198[30]}}, product198});
  assign add_temp_196 = add_signext_392 + add_signext_393;
  assign sum197 = add_temp_196[35:0];

  assign add_signext_394 = sum197;
  assign add_signext_395 = $signed({{5{product199[30]}}, product199});
  assign add_temp_197 = add_signext_394 + add_signext_395;
  assign sum198 = add_temp_197[35:0];

  assign add_signext_396 = sum198;
  assign add_signext_397 = $signed({{5{product200[30]}}, product200});
  assign add_temp_198 = add_signext_396 + add_signext_397;
  assign sum199 = add_temp_198[35:0];

  assign add_signext_398 = sum199;
  assign add_signext_399 = $signed({{5{product201[30]}}, product201});
  assign add_temp_199 = add_signext_398 + add_signext_399;
  assign sum200 = add_temp_199[35:0];

  assign add_signext_400 = sum200;
  assign add_signext_401 = $signed({{5{product202[30]}}, product202});
  assign add_temp_200 = add_signext_400 + add_signext_401;
  assign sum201 = add_temp_200[35:0];

  assign add_signext_402 = sum201;
  assign add_signext_403 = $signed({{5{product203[30]}}, product203});
  assign add_temp_201 = add_signext_402 + add_signext_403;
  assign sum202 = add_temp_201[35:0];

  assign add_signext_404 = sum202;
  assign add_signext_405 = $signed({{5{product204[30]}}, product204});
  assign add_temp_202 = add_signext_404 + add_signext_405;
  assign sum203 = add_temp_202[35:0];

  assign add_signext_406 = sum203;
  assign add_signext_407 = $signed({{5{product205[30]}}, product205});
  assign add_temp_203 = add_signext_406 + add_signext_407;
  assign sum204 = add_temp_203[35:0];

  assign add_signext_408 = sum204;
  assign add_signext_409 = $signed({{5{product206[30]}}, product206});
  assign add_temp_204 = add_signext_408 + add_signext_409;
  assign sum205 = add_temp_204[35:0];

  assign add_signext_410 = sum205;
  assign add_signext_411 = $signed({{5{product207[30]}}, product207});
  assign add_temp_205 = add_signext_410 + add_signext_411;
  assign sum206 = add_temp_205[35:0];

  assign add_signext_412 = sum206;
  assign add_signext_413 = $signed({{5{product208[30]}}, product208});
  assign add_temp_206 = add_signext_412 + add_signext_413;
  assign sum207 = add_temp_206[35:0];

  assign add_signext_414 = sum207;
  assign add_signext_415 = $signed({{5{product209[30]}}, product209});
  assign add_temp_207 = add_signext_414 + add_signext_415;
  assign sum208 = add_temp_207[35:0];

  assign add_signext_416 = sum208;
  assign add_signext_417 = $signed({{5{product210[30]}}, product210});
  assign add_temp_208 = add_signext_416 + add_signext_417;
  assign sum209 = add_temp_208[35:0];

  assign add_signext_418 = sum209;
  assign add_signext_419 = $signed({{5{product211[30]}}, product211});
  assign add_temp_209 = add_signext_418 + add_signext_419;
  assign sum210 = add_temp_209[35:0];

  assign add_signext_420 = sum210;
  assign add_signext_421 = $signed({{5{product212[30]}}, product212});
  assign add_temp_210 = add_signext_420 + add_signext_421;
  assign sum211 = add_temp_210[35:0];

  always @ (posedge clk or posedge reset)
    begin: Output_Register_process
      if (reset == 1'b1) begin
        output_register <= 0;
      end
      else begin
        if (clk_enable == 1'b1) begin
          output_register <= sum211;
        end
      end
    end // Output_Register_process

  // Assignment Statements
  assign filter_out = output_register;
endmodule  // filter1
